netcdf StringAttributes {
  :Conventions = "CF-1.7" ;
}