netcdf nug_atomic_types_enhanced {   // Test
  dimensions:
      dim = 3 ;
  variables:

      char vchar(dim) ;
          vchar:valid_range = "a", "g" ;
      string vstring(dim) ;
          vstring:valid_range = "aaa", "zzzaaaggg" ;

      byte vbyte(dim) ;
          vbyte:valid_range = -5b, 5b ;
      ubyte vubyte(dim) ;
          vubyte:valid_range = 0ub, 6ub ;

      short vshort(dim) ;
          vshort:valid_range = -10s, 10s ;
      ushort vushort(dim) ;
          vushort:valid_range = 0us,  7us;

      int vint(dim) ;
          vint:valid_range = -15, 15 ;
      long vlong(dim) ;
          vlong:valid_range = -20, 20 ;
      uint vuint(dim) ;
          vuint:valid_range = 0u, 15u ;

      int64 vint64(dim) ;
          vint64:valid_range = 0ll, 20ll ;
      uint64 vuint64(dim) ;
          vuint64:valid_range = 0ull, 25ull ;

      float vfloat(dim) ;
          vfloat:valid_range = -25.0f, 25.0f ;
      real vreal(dim) ;
          vreal:valid_range = -30.0f, 30.0f ;

      double vdouble(dim) ;
          vdouble:valid_range = -35.0, 35.0;

  // global attributes
      :title = "test additional atomic data types in enhanced data model" ;

  data:
      vchar   =      "a",    "d",     "g" ;
      vstring = "aaaaaa", "bbbb", "zzaaa" ;

      vbyte   =  -3,  4,  5 ;
      vubyte  =   0,  6,  7 ;

      vshort  =  -4,  9, 10 ;
      vushort =   0, 11, 12 ;

      vint    =  -5, 14, 15 ;
      vlong   =  -6, 19, 20 ;
      vuint   =   0, 21, 22 ;

      vint64  =  -7, 24, 25 ;
      vuint64 =   0, 26, 27 ;

      vfloat  =  -8, 29, 30 ;
      vreal   =  -9, 34, 35 ;

      vdouble = -10, 39, 40 ;
}
