netcdf SpainSoilTemp {
dimensions:
	depth_below_surface_layer = 4 ;
	bounds_dim = 2 ;
	latitude = 16 ;
	time = 9 ;
	longitude = 16 ;
variables:
	double reftime ;
		string reftime:units = "Hour since 2022-09-07T00:00:00Z" ;
		string reftime:standard_name = "forecast_reference_time" ;
		string reftime:long_name = "GRIB reference time" ;
		string reftime:calendar = "proleptic_gregorian" ;
	double depth_below_surface_layer_bounds(depth_below_surface_layer, bounds_dim) ;
		string depth_below_surface_layer_bounds:units = "m" ;
	double depth_below_surface_layer(depth_below_surface_layer) ;
		string depth_below_surface_layer:units = "m" ;
		string depth_below_surface_layer:positive = "down" ;
		string depth_below_surface_layer:bounds = "depth_below_surface_layer_bounds" ;
	float latitude(latitude) ;
		string latitude:units = "degrees_north" ;
		string latitude:standard_name = "latitude" ;
	double time(time) ;
		string time:units = "Hour since 2022-09-07T00:00:00Z" ;
		string time:standard_name = "time" ;
		string time:long_name = "time" ;
		string time:udunits = "Hour since 2022-09-07T00:00:00Z" ;
	float longitude(longitude) ;
		string longitude:units = "degrees_east" ;
		string longitude:standard_name = "longitude" ;
	float Soil_temperature_depth_below_surface_layer(time, depth_below_surface_layer, latitude, longitude) ;
		string Soil_temperature_depth_below_surface_layer:long_name = "Soil temperature @ Depth below land surface layer" ;
		string Soil_temperature_depth_below_surface_layer:units = "K" ;
		string Soil_temperature_depth_below_surface_layer:Grib_Variable_Id = "VAR_2-0-2_L106_layer" ;
		Soil_temperature_depth_below_surface_layer:Grib2_Parameter = 2, 0, 2 ;
		string Soil_temperature_depth_below_surface_layer:Grib2_Parameter_Discipline = "Land surface products" ;
		string Soil_temperature_depth_below_surface_layer:Grib2_Parameter_Category = "Vegetation/Biomass" ;
		string Soil_temperature_depth_below_surface_layer:Grib2_Parameter_Name = "Soil temperature" ;
		Soil_temperature_depth_below_surface_layer:Grib2_Level_Type = 106 ;
		string Soil_temperature_depth_below_surface_layer:Grib2_Level_Desc = "Depth below land surface" ;
		string Soil_temperature_depth_below_surface_layer:Grib2_Generating_Process_Type = "Forecast" ;
		string Soil_temperature_depth_below_surface_layer:Grib2_Statistical_Process_Type = "UnknownStatType--1" ;
		string Soil_temperature_depth_below_surface_layer:coordinates = "reftime time depth_below_surface_layer latitude longitude " ;
		string Soil_temperature_depth_below_surface_layer:grid_mapping = "LatLon_181X360-0p50S-180p00E" ;
	int LatLon_181X360-0p50S-180p00E ;
		string LatLon_181X360-0p50S-180p00E:grid_mapping_name = "latitude_longitude" ;
		LatLon_181X360-0p50S-180p00E:earth_radius = 6371229. ;

// global attributes:
		string :Originating_or_generating_Center = "US National Weather Service, National Centres for Environmental Prediction (NCEP)" ;
		string :Originating_or_generating_Subcenter = "0" ;
		string :GRIB_table_version = "2,1" ;
		string :Type_of_generating_process = "Forecast" ;
		string :Analysis_or_forecast_generating_process_identifier_defined_by_originating_centre = "Analysis from GFS (Global Forecast System)" ;
		string :Conventions = "CF-1.6" ;
		string :history = "Read using CDM IOSP GribCollection v3" ;
		string :featureType = "GRID" ;
		string :History = "Translated to CF-1.0 Conventions by Netcdf-Java CDM (CFGridCoverageWriter)\nOriginal Dataset = GFS_Global_onedeg_20220907_0000.grib2#SRC; Translation Date = 2022-09-08T03:58:21.091Z" ;
		:geospatial_lat_min = 29.5 ;
		:geospatial_lat_max = 45.5 ;
		:geospatial_lon_min = -10.5 ;
		:geospatial_lon_max = 5.5 ;
data:

 reftime = 0 ;

 depth_below_surface_layer_bounds =
  0, 0.100000001490116,
  0.100000001490116, 0.400000005960464,
  0.400000005960464, 1,
  1, 2 ;

 depth_below_surface_layer = 0.0500000007450581, 0.25000000372529, 
    0.700000002980232, 1.5 ;

 latitude = 45, 44, 43, 42, 41, 40, 39, 38, 37, 36, 35, 34, 33, 32, 31, 30 ;

 time = 0, 6, 12, 18, 24, 30, 36, 42, 48 ;

 longitude = 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 
    363, 364, 365 ;

 Soil_temperature_depth_below_surface_layer =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 294.1, 295.4, 295.4, 
    293.6, 290, 290.9, 295.4,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 295, 296, 298.9, 
    296.5, 292, 295.6, 297.6,
  NaNf, 289.3, 288.9, 289.1, 286.1, 286.2, 289.5, 292.7, 292.7, 290.5, 290.8, 
    294.6, 295.2, NaNf, NaNf, NaNf,
  NaNf, NaNf, 288.1, 287, 293, 294.4, 293.5, 289.5, 296.1, 300, 298.4, 295.9, 
    296.4, 298.8, NaNf, NaNf,
  NaNf, NaNf, 289.6, 296, 293.6, 295.1, 292.3, 293.6, 293.5, 297.1, 300.8, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.4, 295.1, 295.5, 295.6, 298.3, 297.5, 295.2, 294.8, 301.8, 
    NaNf, NaNf, NaNf, 300.5, NaNf,
  NaNf, 295.6, 296.1, 296.9, 297.4, 296, 298.7, 298.3, 298.7, 299.4, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.9, 295.7, 298.3, 298.8, 301.8, 298.1, 298.2, 303, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.9, 298.9, 297.9, 298.3, 302.7, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 307.3, 
    304.7, 303.1, 304.2, 302.4,
  NaNf, NaNf, NaNf, NaNf, 298, 299.6, 302.1, 304.7, 301.5, 301.6, 303.4, 
    301.5, 303.2, 303.8, 302.2, 308,
  NaNf, NaNf, NaNf, NaNf, 300.4, 300.7, 301.6, 302.1, 303.4, 302.6, 304.5, 
    303, 301.8, 306, 307.2, 309.9,
  NaNf, NaNf, 298.1, 298.8, 301.7, 298.3, 304.2, 301.1, 302, 302.9, 303.4, 
    305.8, 307, 308.1, 309.1, 310.4,
  NaNf, 299.9, 301.2, 302.3, 295.4, 303.1, 305.9, 308.5, 305.8, 307.8, 306.8, 
    308, 308.7, 309, 309.8, 311.6,
  NaNf, 300.1, 298.1, 305.4, 304.3, 310.1, 310.3, 310.1, 308.6, 308.5, 308.3, 
    309.1, 309.1, 309.6, 310.9, 312.4,
  NaNf, 303.1, 305.4, 310.7, 310.7, 310.5, 312.1, 311.5, 310.2, 309.7, 309.4, 
    309.4, 310.9, 310.8, 310.7, 310.8,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.0925, 292.4925, 
    291.1925, 289.9925, 287.2925, 288.2925, 292.4925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.2925, 292.7925, 
    294.7925, 293.2925, 290.4925, 294.4925, 295.2925,
  NaNf, 289.0925, 288.3925, 288.8925, 286.7925, 287.1925, 288.4925, 290.6925, 
    290.0925, 288.4925, 288.2925, 290.5925, 292.1925, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.5925, 289.7925, 293.9925, 295.9925, 293.9925, 289.2925, 
    295.7925, 298.9925, 298.5925, 295.7925, 295.0925, 295.7925, NaNf, NaNf,
  NaNf, NaNf, 290.5925, 297.0925, 294.3925, 295.9925, 292.3925, 293.7925, 
    293.7925, 296.7925, 299.7925, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.6925, 295.9925, 295.8925, 296.4925, 298.6925, 297.9925, 
    294.9925, 294.9925, 303.8925, NaNf, NaNf, NaNf, 300.8925, NaNf,
  NaNf, 294.4925, 294.9925, 296.7925, 297.5925, 296.2925, 298.6925, 298.5925, 
    298.4925, 299.0925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.2925, 294.4925, 296.0925, 297.3925, 301.0925, 298.4925, 
    298.2925, 302.4925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.5925, 298.2925, 297.4925, 297.8925, 303.9925, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.9925, 
    303.0925, 303.2925, 303.6925, 301.9925,
  NaNf, NaNf, NaNf, NaNf, 299.3925, 298.2925, 302.2925, 304.0925, 303.2925, 
    303.4925, 303.6925, 302.4925, 303.5925, 304.5925, 302.9925, 305.4925,
  NaNf, NaNf, NaNf, NaNf, 301.2925, 302.3925, 302.3925, 302.9925, 304.2925, 
    302.9925, 304.6925, 303.7925, 302.6925, 305.4925, 307.1925, 308.3925,
  NaNf, NaNf, 300.2925, 301.3925, 303.4925, 298.6925, 305.0925, 301.3925, 
    302.1925, 303.0925, 304.6925, 305.6925, 306.6925, 306.8925, 307.8925, 
    309.1925,
  NaNf, 301.7925, 304.3925, 304.2925, 296.4925, 303.2925, 304.6925, 307.5925, 
    305.8925, 307.1925, 306.8925, 307.3925, 307.6925, 307.6925, 308.7925, 
    309.6925,
  NaNf, 299.9925, 299.0925, 305.3925, 304.1925, 308.8925, 309.0925, 308.3925, 
    308.4925, 307.9925, 306.4925, 306.4925, 306.1925, 307.4925, 309.5925, 
    309.9925,
  NaNf, 304.6925, 305.1925, 309.9925, 309.5925, 309.6925, 310.4925, 310.5925, 
    308.3925, 306.8925, 306.8925, 307.0925, 309.9925, 309.4925, 309.5925, 
    307.8925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1792, 290.8192, 
    289.6892, 288.7992, 286.1492, 287.2292, 290.8492,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.3992, 291.2692, 
    292.0592, 290.5892, 289.1792, 293.0292, 293.1192,
  NaNf, 288.6693, 287.9892, 288.3992, 286.0592, 286.5392, 287.3092, 289.3893, 
    288.8092, 287.5592, 287.4292, 289.3593, 290.6592, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1892, 289.5292, 292.5992, 294.7292, 292.1693, 288.4292, 
    294.1992, 296.4292, 296.1792, 294.5992, 293.3992, 293.8692, NaNf, NaNf,
  NaNf, NaNf, 290.1492, 296.5292, 292.8893, 294.6693, 290.6592, 292.3792, 
    292.6492, 295.1192, 298.0392, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.2092, 295.6393, 294.6492, 295.3292, 297.4592, 296.6792, 
    293.0692, 293.8792, 302.8392, NaNf, NaNf, NaNf, 298.4992, NaNf,
  NaNf, 293.2392, 293.5692, 294.9592, 296.7892, 295.0992, 297.7692, 297.2392, 
    296.1492, 297.0892, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6992, 293.7992, 294.5892, 295.5692, 299.1592, 296.6693, 
    296.3593, 299.9193, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.5592, 296.4992, 295.2692, 296.3392, 302.1592, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8492, 
    300.8392, 300.8893, 301.3992, 299.6792,
  NaNf, NaNf, NaNf, NaNf, 298.6192, 296.1992, 300.5192, 301.9592, 301.6292, 
    302.0492, 301.4392, 300.2592, 301.3593, 302.4592, 301.1592, 303.3492,
  NaNf, NaNf, NaNf, NaNf, 300.1292, 302.0992, 300.4392, 301.3893, 302.6693, 
    301.0892, 302.8992, 301.6693, 300.4092, 303.5292, 304.6992, 305.9392,
  NaNf, NaNf, 299.6192, 300.6393, 302.0092, 297.3692, 303.8392, 299.9992, 
    300.6093, 301.3292, 302.6192, 303.6693, 304.4292, 304.6393, 305.5792, 
    306.5592,
  NaNf, 301.2092, 303.9492, 303.2692, 295.7092, 301.8292, 303.0892, 305.7292, 
    303.9792, 305.2792, 304.9992, 305.3792, 305.5992, 305.5792, 306.3593, 
    307.0492,
  NaNf, 298.3192, 297.8893, 303.5692, 302.7492, 307.0592, 307.0492, 306.1792, 
    306.5592, 306.0492, 304.8192, 304.8092, 304.8792, 305.6393, 307.2192, 
    307.4292,
  NaNf, 303.7492, 303.4492, 308.0892, 307.6592, 307.3092, 308.0692, 307.9692, 
    306.6693, 305.6892, 305.6592, 305.7592, 307.5992, 307.1792, 307.1192, 
    305.9292,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.723, 288.573, 
    287.153, 287.343, 284.613, 285.903, 287.833,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.133, 289.513, 
    288.493, 287.023, 287.023, 289.963, 288.923,
  NaNf, 287.793, 287.063, 287.233, 284.533, 284.983, 285.673, 287.743, 
    287.283, 286.413, 286.433, 287.773, 288.463, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.213, 287.483, 288.993, 290.813, 287.623, 286.923, 290.873, 
    292.003, 291.183, 291.893, 289.783, 291.063, NaNf, NaNf,
  NaNf, NaNf, 288.393, 293.513, 288.403, 290.423, 286.893, 289.053, 290.173, 
    292.153, 294.783, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.923, 293.513, 290.633, 291.383, 293.913, 292.433, 289.103, 
    291.043, 301.393, NaNf, NaNf, NaNf, 293.783, NaNf,
  NaNf, 290.613, 290.283, 290.563, 293.203, 291.413, 294.293, 293.773, 
    291.623, 294.243, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.883, 291.883, 291.333, 291.623, 294.063, 292.093, 293.653, 
    296.143, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.323, 292.143, 291.203, 293.833, 299.073, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.283, 
    297.743, 297.843, 298.503, 296.913,
  NaNf, NaNf, NaNf, NaNf, 295.533, 292.363, 297.753, 299.033, 298.313, 
    299.203, 297.993, 297.063, 298.493, 299.573, 298.653, 300.623,
  NaNf, NaNf, NaNf, NaNf, 296.703, 299.973, 297.543, 298.673, 299.833, 
    298.353, 300.173, 299.063, 297.683, 300.723, 301.503, 302.833,
  NaNf, NaNf, 297.103, 298.143, 298.273, 295.373, 301.293, 297.903, 298.333, 
    298.913, 299.983, 300.833, 301.423, 301.643, 302.443, 303.333,
  NaNf, 299.183, 301.683, 300.023, 294.353, 299.703, 300.573, 302.793, 
    301.203, 302.373, 302.093, 302.463, 302.633, 302.653, 303.113, 303.753,
  NaNf, 295.163, 296.313, 301.233, 300.403, 304.053, 303.973, 303.163, 
    304.013, 303.113, 302.243, 302.313, 303.023, 302.953, 303.933, 304.133,
  NaNf, 301.543, 300.953, 304.983, 304.543, 304.103, 304.843, 304.683, 
    304.143, 303.863, 303.783, 303.803, 304.283, 303.963, 303.883, 303.463,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4925, 294.0925, 
    293.8925, 292.3925, 288.9925, 289.8925, 293.6925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.5925, 294.3925, 
    296.1925, 294.2925, 290.7925, 293.9925, 295.8925,
  NaNf, 288.7925, 287.9925, 287.7925, 284.4925, 284.7925, 287.6925, 290.9925, 
    291.0925, 289.1925, 289.3925, 293.0925, 293.3925, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.0925, 285.5925, 290.3925, 290.6925, 289.8925, 287.4925, 
    292.1925, 296.0925, 295.4925, 293.4925, 293.7925, 296.6925, NaNf, NaNf,
  NaNf, NaNf, 288.2925, 292.1925, 290.4925, 291.1925, 288.8925, 290.5925, 
    289.9925, 293.3925, 297.4925, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.5925, 291.5925, 292.5925, 292.4925, 294.2925, 293.2925, 
    291.7925, 290.9925, 299.6925, NaNf, NaNf, NaNf, 298.1925, NaNf,
  NaNf, 293.2925, 293.6925, 294.0925, 293.8925, 293.1925, 294.4925, 294.1925, 
    295.1925, 295.7925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.2925, 293.0925, 295.0925, 295.6925, 297.8925, 294.4925, 
    293.7925, 299.1925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 296.4925, 295.1925, 293.9925, 294.4925, 298.7925, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 303.3925, 
    301.1925, 300.1925, 300.6925, 300.1925,
  NaNf, NaNf, NaNf, NaNf, 295.0925, 295.9925, 297.6925, 300.7925, 299.0925, 
    299.6925, 299.8925, 298.4925, 299.5925, 300.3925, 299.4925, 304.4925,
  NaNf, NaNf, NaNf, NaNf, 296.3925, 297.1925, 297.1925, 298.3925, 300.5925, 
    299.0925, 300.3925, 299.7925, 297.9925, 301.4925, 303.6925, 306.0925,
  NaNf, NaNf, 294.8925, 294.7925, 297.3925, 293.8925, 299.3925, 296.8925, 
    298.5925, 298.1925, 299.4925, 301.9925, 303.2925, 303.8925, 304.5925, 
    306.4925,
  NaNf, 295.7925, 296.6925, 297.8925, 291.2925, 298.2925, 301.1925, 304.6925, 
    301.6925, 303.2925, 302.8925, 303.8925, 304.9925, 305.0925, 305.6925, 
    307.5925,
  NaNf, 295.6925, 293.0925, 300.0925, 298.9925, 304.7925, 305.9925, 305.2925, 
    304.4925, 304.7925, 305.2925, 306.0925, 306.2925, 306.1925, 306.8925, 
    308.3925,
  NaNf, 297.6925, 299.8925, 305.3925, 305.4925, 305.7925, 307.1925, 306.7925, 
    306.4925, 306.4925, 306.4925, 306.5925, 307.4925, 306.8925, 306.7925, 
    307.5925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.0162, 292.5063, 
    291.2162, 289.9763, 287.2362, 288.2662, 292.5063,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.2762, 292.7863, 
    294.8163, 293.2963, 290.5363, 294.4662, 295.3463,
  NaNf, 289.0963, 288.4362, 288.8662, 286.6862, 287.1762, 288.4463, 290.6363, 
    290.0463, 288.4562, 288.2863, 290.6462, 292.1963, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.5862, 289.6063, 293.8362, 295.7263, 293.8362, 289.2263, 
    295.7263, 298.8463, 298.4662, 295.6663, 295.0363, 295.8062, NaNf, NaNf,
  NaNf, NaNf, 290.6063, 296.9163, 294.2963, 295.8563, 292.2863, 293.6562, 
    293.6263, 296.6862, 299.6562, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.5963, 295.9163, 295.8463, 296.3863, 298.5663, 297.7963, 
    294.8463, 294.8662, 303.2662, NaNf, NaNf, NaNf, 300.7563, NaNf,
  NaNf, 294.4862, 295.0063, 296.7462, 297.4862, 296.1862, 298.4862, 298.4362, 
    298.3563, 298.9362, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.2062, 294.4662, 296.0562, 297.3362, 301.0162, 298.3662, 
    298.0862, 302.3163, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.4562, 298.2362, 297.3362, 297.7662, 303.8062, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.8362, 
    303.0063, 303.0663, 303.5862, 301.8962,
  NaNf, NaNf, NaNf, NaNf, 299.2162, 298.2563, 302.0463, 303.8863, 303.0763, 
    303.1862, 303.4763, 302.3163, 303.3662, 304.3563, 302.8463, 305.3763,
  NaNf, NaNf, NaNf, NaNf, 301.0862, 301.9362, 302.0663, 302.7662, 304.1063, 
    302.7062, 304.5162, 303.5763, 302.4262, 305.3863, 307.0262, 308.3062,
  NaNf, NaNf, 299.9763, 301.1562, 303.1562, 298.4763, 304.9262, 301.1462, 
    301.9962, 302.8263, 304.3662, 305.4962, 306.4763, 306.7462, 307.7462, 
    309.0463,
  NaNf, 301.6562, 304.1562, 304.0063, 296.3062, 303.1562, 304.5562, 307.4763, 
    305.7263, 307.0463, 306.7563, 307.2563, 307.5562, 307.5763, 308.6663, 
    309.5562,
  NaNf, 299.8463, 298.7863, 305.1862, 304.0763, 308.7762, 308.9962, 308.2263, 
    308.2563, 307.8163, 306.4362, 306.4562, 306.1363, 307.4562, 309.5063, 
    309.9562,
  NaNf, 304.3662, 305.0363, 309.8662, 309.4463, 309.5162, 310.3463, 310.4062, 
    308.3163, 306.8763, 306.8763, 307.0562, 309.8863, 309.3962, 309.3962, 
    307.7662,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1885, 290.8385, 
    289.6885, 288.7985, 286.1485, 287.2285, 290.8585,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4085, 291.2785, 
    292.0685, 290.5985, 289.1885, 293.0385, 293.1285,
  NaNf, 288.6685, 287.9885, 288.3985, 286.0585, 286.5385, 287.3185, 289.3885, 
    288.8185, 287.5685, 287.4385, 289.3685, 290.6585, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1785, 289.5085, 292.5885, 294.7185, 292.1685, 288.4285, 
    294.1985, 296.4285, 296.1785, 294.5985, 293.3985, 293.8785, NaNf, NaNf,
  NaNf, NaNf, 290.1485, 296.5085, 292.8785, 294.6585, 290.6485, 292.3685, 
    292.6485, 295.1185, 298.0385, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.2085, 295.6285, 294.6385, 295.3185, 297.4485, 296.6585, 
    293.0685, 293.8785, 302.8385, NaNf, NaNf, NaNf, 298.5085, NaNf,
  NaNf, 293.2385, 293.5685, 294.9485, 296.7685, 295.0885, 297.7485, 297.2385, 
    296.1385, 297.0985, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6885, 293.7885, 294.5785, 295.5685, 299.1485, 296.6585, 
    296.3685, 299.9185, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.5385, 296.4885, 295.2685, 296.3385, 302.1585, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8585, 
    300.8485, 300.8985, 301.4085, 299.6885,
  NaNf, NaNf, NaNf, NaNf, 298.5985, 296.1885, 300.5185, 301.9685, 301.6185, 
    302.0485, 301.4385, 300.2585, 301.3685, 302.4685, 301.1685, 303.3585,
  NaNf, NaNf, NaNf, NaNf, 300.1085, 302.0685, 300.4485, 301.3885, 302.6685, 
    301.0885, 302.9085, 301.6785, 300.4285, 303.5385, 304.7085, 305.9585,
  NaNf, NaNf, 299.5985, 300.6185, 301.9985, 297.3785, 303.8285, 299.9985, 
    300.6085, 301.3385, 302.6285, 303.6785, 304.4385, 304.6485, 305.5885, 
    306.5685,
  NaNf, 301.1985, 303.9285, 303.2585, 295.7085, 301.8385, 303.0985, 305.7285, 
    303.9885, 305.2885, 304.9985, 305.3885, 305.5985, 305.5885, 306.3685, 
    307.0685,
  NaNf, 298.3185, 297.8885, 303.5785, 302.7485, 307.0585, 307.0485, 306.1885, 
    306.5685, 306.0585, 304.8185, 304.8085, 304.8885, 305.6485, 307.2285, 
    307.4385,
  NaNf, 303.7385, 303.4585, 308.0885, 307.6685, 307.3185, 308.0785, 307.9785, 
    306.6785, 305.6885, 305.6685, 305.7685, 307.6085, 307.1885, 307.1285, 
    305.9385,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.723, 288.583, 
    287.163, 287.353, 284.623, 285.913, 287.843,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.143, 289.523, 
    288.503, 287.033, 287.033, 289.973, 288.933,
  NaNf, 287.793, 287.073, 287.243, 284.543, 284.993, 285.683, 287.753, 
    287.293, 286.423, 286.443, 287.783, 288.473, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.213, 287.493, 289.003, 290.833, 287.633, 286.933, 290.883, 
    292.013, 291.193, 291.903, 289.793, 291.073, NaNf, NaNf,
  NaNf, NaNf, 288.403, 293.513, 288.413, 290.433, 286.903, 289.063, 290.183, 
    292.173, 294.793, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.923, 293.523, 290.643, 291.393, 293.923, 292.443, 289.113, 
    291.053, 301.393, NaNf, NaNf, NaNf, 293.793, NaNf,
  NaNf, 290.623, 290.293, 290.563, 293.213, 291.423, 294.303, 293.783, 
    291.633, 294.263, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.883, 291.893, 291.343, 291.633, 294.073, 292.103, 293.663, 
    296.153, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.333, 292.153, 291.213, 293.843, 299.093, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.303, 
    297.763, 297.853, 298.513, 296.923,
  NaNf, NaNf, NaNf, NaNf, 295.543, 292.383, 297.763, 299.043, 298.333, 
    299.213, 298.013, 297.083, 298.503, 299.593, 298.663, 300.633,
  NaNf, NaNf, NaNf, NaNf, 296.713, 299.973, 297.553, 298.683, 299.843, 
    298.363, 300.183, 299.083, 297.703, 300.743, 301.523, 302.843,
  NaNf, NaNf, 297.103, 298.153, 298.283, 295.383, 301.303, 297.913, 298.343, 
    298.923, 299.993, 300.853, 301.433, 301.663, 302.453, 303.343,
  NaNf, 299.183, 301.693, 300.033, 294.363, 299.713, 300.583, 302.803, 
    301.213, 302.383, 302.113, 302.483, 302.643, 302.663, 303.133, 303.773,
  NaNf, 295.173, 296.323, 301.243, 300.413, 304.063, 303.983, 303.173, 
    304.033, 303.123, 302.253, 302.323, 303.033, 302.963, 303.953, 304.153,
  NaNf, 301.543, 300.963, 304.993, 304.553, 304.113, 304.853, 304.693, 
    304.163, 303.873, 303.793, 303.813, 304.293, 303.973, 303.903, 303.473,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.6, 294.8, 294.1, 
    292.7, 289.6, 290.8, 295.2,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 294.5, 295.1, 298.2, 
    295.3, 292.2, 295.6, 298,
  NaNf, 289.3, 288.3, 288.4, 285.4, 285.9, 288.6, 291.9, 291.8, 289.9, 290.3, 
    293.5, 294.4, NaNf, NaNf, NaNf,
  NaNf, NaNf, 288, 286.5, 292.4, 294.9, 292.8, 288.3, 294.9, 299.1, 299.3, 
    297, 297, 299.1, NaNf, NaNf,
  NaNf, NaNf, 288.8, 294.6, 292, 294.8, 290.9, 292.5, 291.9, 296.5, 301.8, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 290.4, 293.7, 293.3, 293.7, 297.5, 298, 295.6, 296.4, 307.6, 
    NaNf, NaNf, NaNf, 303, NaNf,
  NaNf, 295.4, 295.1, 295.9, 296.5, 295, 298.7, 299, 299.3, 301.3, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.5, 294.4, 296.7, 298.1, 301.9, 298.8, 300.8, 305.2, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 301.3, 299.2, 298.6, 300.2, 308, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 310.2, 
    305.7, 307.6, 307.1, 306.6,
  NaNf, NaNf, NaNf, NaNf, 300.1, 299.6, 306, 309, 307, 308.4, 306.4, 303.9, 
    306.5, 308.4, 306, 310.2,
  NaNf, NaNf, NaNf, NaNf, 302.6, 303.3, 304.9, 306.6, 307.3, 303.3, 307.1, 
    307.2, 305.5, 308.7, 311.4, 313.7,
  NaNf, NaNf, 301.2, 301, 305.4, 301, 307.3, 303.6, 304.5, 303.3, 304.9, 
    308.6, 308.4, 309.8, 311.6, 314,
  NaNf, 301.5, 304.5, 304.5, 298.4, 306.2, 307.4, 309.9, 307.6, 309.1, 309, 
    310.3, 310.2, 311.3, 312.3, 314.3,
  NaNf, 301.6, 301.9, 308.6, 306, 312.1, 311.8, 309.5, 311.3, 310.1, 309.4, 
    309.7, 309.8, 311.2, 313.1, 314.6,
  NaNf, 306.3, 307.7, 312.3, 312.4, 312.5, 313.2, 313, 310.9, 309.9, 310.2, 
    310.3, 312.9, 312.7, 313, 312.3,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.9, 292.5, 291.2, 
    290, 287.2, 288.3, 292.5,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.2, 292.8, 294.8, 
    293.2, 290.5, 294.4, 295.3,
  NaNf, 289.1, 288.4, 288.8, 286.6, 287.1, 288.4, 290.6, 290, 288.4, 288.3, 
    290.6, 292.2, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.5, 289.5, 293.7, 295.5, 293.6, 289.1, 295.5, 298.6, 298.3, 
    295.6, 294.9, 295.8, NaNf, NaNf,
  NaNf, NaNf, 290.5, 296.7, 294.2, 295.7, 292.2, 293.5, 293.5, 296.5, 299.6, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.5, 295.7, 295.7, 296.2, 298.4, 297.6, 294.8, 294.7, 303.2, 
    NaNf, NaNf, NaNf, 300.6, NaNf,
  NaNf, 294.4, 294.9, 296.7, 297.4, 296.1, 298.3, 298.3, 298.2, 298.8, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297, 294.5, 296, 297.3, 300.9, 298.3, 297.9, 302.2, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.4, 298.1, 297.2, 297.7, 303.7, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.7, 
    302.9, 303, 303.4, 301.8,
  NaNf, NaNf, NaNf, NaNf, 299.1, 298.2, 301.9, 303.8, 302.9, 303.1, 303.3, 
    302.2, 303.2, 304.2, 302.7, 305.4,
  NaNf, NaNf, NaNf, NaNf, 300.9, 301.7, 301.9, 302.6, 304, 302.5, 304.3, 
    303.4, 302.3, 305.3, 306.9, 308.2,
  NaNf, NaNf, 299.8, 301, 302.9, 298.3, 304.7, 301, 301.9, 302.6, 304.2, 
    305.4, 306.4, 306.7, 307.7, 309,
  NaNf, 301.5, 303.9, 303.7, 296.1, 303, 304.4, 307.3, 305.6, 306.9, 306.6, 
    307.1, 307.4, 307.5, 308.6, 309.5,
  NaNf, 299.7, 298.6, 305, 303.9, 308.6, 308.8, 308.1, 308.1, 307.7, 306.3, 
    306.4, 306.1, 307.4, 309.4, 309.9,
  NaNf, 304.1, 304.9, 309.7, 309.3, 309.3, 310.1, 310.2, 308.2, 306.8, 306.8, 
    307, 309.7, 309.3, 309.3, 307.7,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1892, 290.8392, 
    289.6992, 288.8092, 286.1592, 287.2392, 290.8692,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4092, 291.2892, 
    292.0792, 290.6093, 289.1892, 293.0392, 293.1393,
  NaNf, 288.6693, 287.9892, 288.3893, 286.0492, 286.5292, 287.3192, 289.3992, 
    288.8292, 287.5692, 287.4492, 289.3792, 290.6693, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1592, 289.4892, 292.5792, 294.6892, 292.1492, 288.4292, 
    294.1892, 296.4292, 296.1792, 294.5992, 293.3992, 293.8792, NaNf, NaNf,
  NaNf, NaNf, 290.1393, 296.4792, 292.8593, 294.6393, 290.6492, 292.3593, 
    292.6393, 295.1192, 298.0392, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1992, 295.6093, 294.6192, 295.2992, 297.4292, 296.6393, 
    293.0592, 293.8692, 302.8092, NaNf, NaNf, NaNf, 298.5192, NaNf,
  NaNf, 293.2392, 293.5692, 294.9392, 296.7492, 295.0692, 297.7192, 297.2092, 
    296.1393, 297.0992, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6693, 293.7892, 294.5692, 295.5592, 299.1393, 296.6492, 
    296.3692, 299.9292, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.5292, 296.4792, 295.2692, 296.3392, 302.1492, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8492, 
    300.8593, 300.9092, 301.4193, 299.6992,
  NaNf, NaNf, NaNf, NaNf, 298.5792, 296.1892, 300.5192, 301.9692, 301.6093, 
    302.0292, 301.4392, 300.2692, 301.3692, 302.4692, 301.1693, 303.3593,
  NaNf, NaNf, NaNf, NaNf, 300.0892, 302.0192, 300.4392, 301.3792, 302.6592, 
    301.0892, 302.8992, 301.6792, 300.4292, 303.5392, 304.7192, 305.9692,
  NaNf, NaNf, 299.5792, 300.5992, 301.9692, 297.3692, 303.8192, 299.9992, 
    300.6093, 301.3292, 302.6292, 303.6792, 304.4492, 304.6492, 305.5992, 
    306.5792,
  NaNf, 301.1792, 303.8992, 303.2292, 295.6992, 301.8392, 303.0892, 305.7292, 
    303.9892, 305.2892, 304.9992, 305.3893, 305.6093, 305.5892, 306.3792, 
    307.0792,
  NaNf, 298.3092, 297.8893, 303.5792, 302.7492, 307.0592, 307.0592, 306.1892, 
    306.5692, 306.0592, 304.8192, 304.8192, 304.8893, 305.6492, 307.2392, 
    307.4592,
  NaNf, 303.7192, 303.4592, 308.0892, 307.6592, 307.3292, 308.0892, 307.9892, 
    306.6792, 305.6992, 305.6693, 305.7692, 307.6093, 307.1892, 307.1292, 
    305.9492,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.7337, 288.5937, 
    287.1637, 287.3537, 284.6237, 285.9237, 287.8537,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.1437, 289.5337, 
    288.5137, 287.0437, 287.0437, 289.9837, 288.9437,
  NaNf, 287.8037, 287.0737, 287.2537, 284.5537, 285.0037, 285.6837, 287.7537, 
    287.3037, 286.4237, 286.4537, 287.7837, 288.4837, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.2237, 287.5037, 289.0137, 290.8437, 287.6437, 286.9437, 
    290.9037, 292.0237, 291.2037, 291.9137, 289.8037, 291.0837, NaNf, NaNf,
  NaNf, NaNf, 288.4037, 293.5237, 288.4337, 290.4437, 286.9137, 289.0737, 
    290.1837, 292.1837, 294.8037, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.9337, 293.5137, 290.6537, 291.4037, 293.9337, 292.4537, 
    289.1237, 291.0637, 301.3937, NaNf, NaNf, NaNf, 293.8037, NaNf,
  NaNf, 290.6237, 290.3037, 290.5737, 293.2237, 291.4337, 294.3137, 293.7937, 
    291.6437, 294.2737, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.8937, 291.9037, 291.3537, 291.6437, 294.0837, 292.1137, 
    293.6737, 296.1637, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.3437, 292.1637, 291.2237, 293.8537, 299.1037, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.3137, 
    297.7737, 297.8637, 298.5237, 296.9337,
  NaNf, NaNf, NaNf, NaNf, 295.5537, 292.3937, 297.7737, 299.0537, 298.3437, 
    299.2237, 298.0337, 297.0937, 298.5237, 299.6037, 298.6737, 300.6437,
  NaNf, NaNf, NaNf, NaNf, 296.7237, 299.9737, 297.5737, 298.6937, 299.8537, 
    298.3737, 300.1937, 299.0937, 297.7137, 300.7537, 301.5337, 302.8637,
  NaNf, NaNf, 297.1137, 298.1637, 298.2937, 295.3937, 301.3137, 297.9237, 
    298.3537, 298.9337, 300.0037, 300.8637, 301.4437, 301.6737, 302.4737, 
    303.3537,
  NaNf, 299.1937, 301.6937, 300.0437, 294.3737, 299.7237, 300.5937, 302.8237, 
    301.2237, 302.3937, 302.1237, 302.4937, 302.6637, 302.6837, 303.1437, 
    303.7837,
  NaNf, 295.1837, 296.3237, 301.2437, 300.4237, 304.0737, 303.9937, 303.1837, 
    304.0437, 303.1337, 302.2737, 302.3337, 303.0437, 302.9737, 303.9637, 
    304.1637,
  NaNf, 301.5537, 300.9737, 305.0037, 304.5637, 304.1237, 304.8737, 304.7137, 
    304.1737, 303.8837, 303.7937, 303.8237, 304.3137, 303.9837, 303.9137, 
    303.4837,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 294.3925, 295.6925, 
    294.9925, 293.1925, 290.2925, 291.3925, 296.2925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 295.2925, 296.2925, 
    299.6925, 296.8925, 292.8925, 296.4925, 299.1925,
  NaNf, 290.1925, 289.1925, 289.2925, 286.1925, 286.5925, 289.5925, 293.0925, 
    292.6925, 290.5925, 290.6925, 294.2925, 295.6925, NaNf, NaNf, NaNf,
  NaNf, NaNf, 288.9925, 287.8925, 294.3925, 297.7925, 294.7925, 289.2925, 
    296.6925, 301.6925, 301.1925, 298.5925, 299.2925, 300.4925, NaNf, NaNf,
  NaNf, NaNf, 289.7925, 297.8925, 294.3925, 296.8925, 291.9925, 294.1925, 
    293.7925, 298.7925, 304.3925, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.7925, 296.6925, 295.4925, 295.9925, 299.1925, 299.5925, 
    297.2925, 298.4925, 307.2925, NaNf, NaNf, NaNf, 304.3925, NaNf,
  NaNf, 297.4925, 297.1925, 298.2925, 299.4925, 297.5925, 301.9925, 302.0925, 
    302.1925, 304.0925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 301.1925, 296.8925, 299.3925, 300.5925, 305.1925, 302.0925, 
    303.8925, 308.9925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 304.1925, 302.4925, 302.1925, 303.7925, 310.6925, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 313.4925, 
    308.1925, 309.6925, 309.5925, 308.4925,
  NaNf, NaNf, NaNf, NaNf, 302.7925, 303.3925, 308.7925, 310.7925, 308.8925, 
    307.8925, 310.1925, 306.6925, 309.5925, 309.9925, 308.3925, 312.4925,
  NaNf, NaNf, NaNf, NaNf, 306.3925, 305.8925, 308.8925, 309.8925, 309.5925, 
    306.7925, 310.1925, 308.3925, 307.6925, 310.9925, 313.5925, 316.1925,
  NaNf, NaNf, 305.0925, 305.6925, 308.6925, 304.5925, 311.8925, 306.0925, 
    307.6925, 306.9925, 308.7925, 309.7925, 311.6925, 311.0925, 313.0925, 
    316.6925,
  NaNf, 307.0925, 310.1925, 310.1925, 301.9925, 310.3925, 310.9925, 313.6925, 
    310.1925, 310.8925, 311.6925, 312.5925, 312.9925, 313.2925, 315.0925, 
    316.7925,
  NaNf, 306.0925, 307.0925, 312.9925, 310.2925, 316.8925, 315.5925, 313.0925, 
    314.7925, 312.7925, 311.7925, 311.9925, 312.5925, 313.7925, 315.8925, 
    316.6925,
  NaNf, 311.8925, 312.5925, 317.2925, 317.6925, 316.9925, 317.8925, 317.6925, 
    314.2925, 312.8925, 313.1925, 313.2925, 315.8925, 315.4925, 315.7925, 
    314.6925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.9, 292.5, 291.2, 
    290, 287.2, 288.3, 292.6,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.3, 292.8, 294.8, 
    293.3, 290.5, 294.4, 295.4,
  NaNf, 289.1, 288.4, 288.8, 286.6, 287.1, 288.4, 290.6, 290, 288.4, 288.3, 
    290.7, 292.2, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.4, 289.4, 293.7, 295.6, 293.6, 289.1, 295.5, 298.7, 298.4, 
    295.7, 295, 295.8, NaNf, NaNf,
  NaNf, NaNf, 290.5, 296.7, 294.1, 295.7, 292.1, 293.5, 293.5, 296.6, 299.8, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.5, 295.8, 295.6, 296.1, 298.4, 297.7, 294.8, 294.9, 304.1, 
    NaNf, NaNf, NaNf, 300.8, NaNf,
  NaNf, 294.5, 294.9, 296.7, 297.4, 296.1, 298.5, 298.4, 298.3, 299, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.2, 294.5, 296, 297.3, 301, 298.3, 298.2, 302.4, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.6, 298.2, 297.3, 297.8, 304, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.9, 
    303, 303.2, 303.7, 302,
  NaNf, NaNf, NaNf, NaNf, 299.2, 298.2, 302.3, 304.1, 303.3, 303.5, 303.6, 
    302.3, 303.5, 304.5, 303, 305.5,
  NaNf, NaNf, NaNf, NaNf, 301.2, 302.2, 302.2, 303, 304.3, 302.7, 304.6, 
    303.7, 302.5, 305.4, 307.2, 308.5,
  NaNf, NaNf, 300.1, 301.1, 303.3, 298.7, 305, 301.3, 302.1, 302.8, 304.4, 
    305.5, 306.5, 306.8, 307.8, 309.2,
  NaNf, 301.6, 304.1, 304, 296.5, 303.2, 304.6, 307.6, 305.7, 307, 306.8, 
    307.3, 307.6, 307.6, 308.7, 309.7,
  NaNf, 299.9, 299, 305.3, 304.1, 309, 309.2, 308.2, 308.4, 307.8, 306.4, 
    306.5, 306.2, 307.5, 309.6, 310.1,
  NaNf, 304.5, 305.1, 309.9, 309.5, 309.7, 310.5, 310.4, 308.3, 306.9, 306.9, 
    307.1, 309.9, 309.5, 309.5, 307.8,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1785, 290.8485, 
    289.6985, 288.8185, 286.1685, 287.2485, 290.8785,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4185, 291.2985, 
    292.0985, 290.6185, 289.1985, 293.0385, 293.1485,
  NaNf, 288.6685, 287.9885, 288.3885, 286.0485, 286.5285, 287.3185, 289.3985, 
    288.8385, 287.5685, 287.4485, 289.3885, 290.6785, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1485, 289.4685, 292.5685, 294.6685, 292.1485, 288.4185, 
    294.1885, 296.4285, 296.1685, 294.5885, 293.3985, 293.8985, NaNf, NaNf,
  NaNf, NaNf, 290.1285, 296.4485, 292.8485, 294.6285, 290.6385, 292.3485, 
    292.6285, 295.1185, 298.0385, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1885, 295.5785, 294.6085, 295.2785, 297.4085, 296.6185, 
    293.0585, 293.8585, 302.8185, NaNf, NaNf, NaNf, 298.5285, NaNf,
  NaNf, 293.2285, 293.5585, 294.9385, 296.7285, 295.0585, 297.6985, 297.1985, 
    296.1385, 297.0985, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6485, 293.7785, 294.5685, 295.5585, 299.1185, 296.6385, 
    296.3685, 299.9285, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.5085, 296.4685, 295.2685, 296.3385, 302.1485, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8485, 
    300.8585, 300.9185, 301.4285, 299.7085,
  NaNf, NaNf, NaNf, NaNf, 298.5685, 296.1885, 300.5185, 301.9785, 301.5985, 
    302.0185, 301.4385, 300.2685, 301.3785, 302.4785, 301.1785, 303.3685,
  NaNf, NaNf, NaNf, NaNf, 300.0785, 301.9785, 300.4385, 301.3785, 302.6585, 
    301.0885, 302.8985, 301.6885, 300.4385, 303.5485, 304.7285, 305.9785,
  NaNf, NaNf, 299.5585, 300.5785, 301.9485, 297.3785, 303.8185, 299.9985, 
    300.6085, 301.3285, 302.6285, 303.6785, 304.4485, 304.6585, 305.6085, 
    306.5985,
  NaNf, 301.1685, 303.8785, 303.2085, 295.6985, 301.8385, 303.0885, 305.7285, 
    303.9885, 305.2885, 305.0085, 305.3885, 305.6085, 305.5985, 306.3885, 
    307.0885,
  NaNf, 298.3085, 297.8885, 303.5785, 302.7385, 307.0585, 307.0585, 306.1985, 
    306.5785, 306.0585, 304.8285, 304.8185, 304.8985, 305.6585, 307.2385, 
    307.4685,
  NaNf, 303.6985, 303.4585, 308.0885, 307.6585, 307.3285, 308.0985, 307.9985, 
    306.6885, 305.6985, 305.6685, 305.7785, 307.6185, 307.1985, 307.1385, 
    305.9685,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.743, 288.603, 
    287.183, 287.373, 284.643, 285.923, 287.863,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.153, 289.543, 
    288.523, 287.053, 287.053, 289.993, 288.953,
  NaNf, 287.803, 287.083, 287.263, 284.553, 285.013, 285.693, 287.773, 
    287.313, 286.433, 286.463, 287.793, 288.493, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.233, 287.513, 289.023, 290.853, 287.663, 286.943, 290.913, 
    292.033, 291.213, 291.923, 289.813, 291.093, NaNf, NaNf,
  NaNf, NaNf, 288.413, 293.533, 288.443, 290.453, 286.923, 289.083, 290.203, 
    292.193, 294.813, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.933, 293.533, 290.663, 291.413, 293.943, 292.473, 289.143, 
    291.073, 301.393, NaNf, NaNf, NaNf, 293.813, NaNf,
  NaNf, 290.633, 290.303, 290.583, 293.233, 291.443, 294.323, 293.803, 
    291.653, 294.283, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.903, 291.913, 291.363, 291.653, 294.103, 292.123, 293.683, 
    296.183, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.353, 292.173, 291.233, 293.863, 299.113, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.333, 
    297.793, 297.883, 298.543, 296.953,
  NaNf, NaNf, NaNf, NaNf, 295.563, 292.403, 297.783, 299.073, 298.353, 
    299.243, 298.043, 297.113, 298.533, 299.613, 298.683, 300.663,
  NaNf, NaNf, NaNf, NaNf, 296.733, 299.973, 297.583, 298.703, 299.863, 
    298.393, 300.203, 299.103, 297.723, 300.763, 301.543, 302.873,
  NaNf, NaNf, 297.123, 298.173, 298.303, 295.403, 301.323, 297.933, 298.363, 
    298.953, 300.013, 300.873, 301.463, 301.683, 302.483, 303.373,
  NaNf, 299.203, 301.703, 300.053, 294.373, 299.733, 300.603, 302.833, 
    301.243, 302.413, 302.133, 302.503, 302.673, 302.693, 303.153, 303.793,
  NaNf, 295.193, 296.333, 301.253, 300.433, 304.083, 304.013, 303.203, 
    304.063, 303.153, 302.283, 302.343, 303.053, 302.983, 303.983, 304.183,
  NaNf, 301.563, 300.983, 305.013, 304.573, 304.143, 304.883, 304.723, 
    304.183, 303.893, 303.813, 303.833, 304.323, 304.003, 303.933, 303.503,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.2, 293.9, 293.5, 
    292, 289.1, 290.2, 294.9,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.6, 294.6, 296.6, 
    294.8, 291.7, 295, 297.1,
  NaNf, 289.7, 288.7, 288.6, 285.1, 285, 288.1, 291.1, 291.3, 289.2, 288.9, 
    292.7, 293.9, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.9, 286.5, 292.2, 293.6, 291.9, 287.9, 293.1, 297.5, 297.8, 
    295.6, 296.7, 298.9, NaNf, NaNf,
  NaNf, NaNf, 289, 295.1, 292.3, 293.4, 289.7, 291.6, 290.8, 294.8, 300, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 290.7, 294.5, 294.2, 294.3, 295.9, 295.3, 294.1, 294.4, 302.2, 
    NaNf, NaNf, NaNf, 301.1, NaNf,
  NaNf, 295.2, 295.6, 296.4, 297, 295.5, 297.9, 297.6, 299, 299.7, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6, 295.4, 297.2, 297.9, 300.8, 297.8, 298.1, 303.8, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.5, 298.4, 297.8, 299, 303.5, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.6, 
    302.8, 303.8, 304.5, 303.8,
  NaNf, NaNf, NaNf, NaNf, 298.2, 299.3, 301.7, 304.2, 302.6, 301.4, 303.6, 
    301.7, 303.8, 304.6, 303.2, 308.2,
  NaNf, NaNf, NaNf, NaNf, 300.4, 300.4, 302, 302.1, 302.7, 301.8, 304.2, 
    302.6, 302.2, 304.9, 307.5, 310.7,
  NaNf, NaNf, 299.1, 299.6, 302, 297.8, 304.7, 300.1, 301.9, 301.9, 302.8, 
    304.8, 306.5, 306.1, 308.8, 311.4,
  NaNf, 301.2, 302.4, 303.8, 295.7, 303.3, 305.1, 307.3, 304.7, 305.9, 307.3, 
    307.8, 308.7, 308.4, 310.2, 311.3,
  NaNf, 300, 298.6, 305.2, 303.6, 310, 309, 307.6, 308.3, 308.2, 308.2, 
    308.1, 309, 309.3, 310.6, 311.3,
  NaNf, 303.4, 305, 310.7, 310.9, 310.6, 311, 311.1, 310, 309.4, 309.5, 
    310.1, 311.3, 310.5, 310.8, 310.2,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.9, 292.5, 291.2, 
    290, 287.2, 288.3, 292.6,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.2, 292.8, 294.9, 
    293.3, 290.5, 294.4, 295.4,
  NaNf, 289.1, 288.4, 288.8, 286.6, 287.1, 288.4, 290.6, 290, 288.4, 288.3, 
    290.7, 292.2, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.4, 289.3, 293.7, 295.5, 293.6, 289.1, 295.5, 298.7, 298.4, 
    295.7, 295.1, 295.9, NaNf, NaNf,
  NaNf, NaNf, 290.5, 296.7, 294.1, 295.6, 292.1, 293.4, 293.4, 296.5, 299.8, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.5, 295.8, 295.6, 296.1, 298.4, 297.6, 294.8, 294.9, 304, 
    NaNf, NaNf, NaNf, 300.8, NaNf,
  NaNf, 294.5, 294.9, 296.6, 297.4, 296.1, 298.5, 298.4, 298.4, 299.1, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.3, 294.5, 296.1, 297.3, 301, 298.4, 298.3, 302.5, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.6, 298.3, 297.4, 297.9, 304.1, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 307, 303, 
    303.3, 303.7, 302.1,
  NaNf, NaNf, NaNf, NaNf, 299.2, 298.3, 302.3, 304.2, 303.3, 303.5, 303.7, 
    302.3, 303.6, 304.6, 303, 305.6,
  NaNf, NaNf, NaNf, NaNf, 301.2, 302.2, 302.3, 303, 304.3, 302.7, 304.7, 
    303.7, 302.5, 305.5, 307.2, 308.6,
  NaNf, NaNf, 300.1, 301.1, 303.3, 298.8, 305.1, 301.3, 302.2, 302.8, 304.4, 
    305.5, 306.5, 306.7, 307.8, 309.3,
  NaNf, 301.7, 304.2, 304.2, 296.6, 303.3, 304.7, 307.6, 305.7, 307, 306.8, 
    307.4, 307.6, 307.6, 308.8, 309.8,
  NaNf, 299.9, 299.1, 305.4, 304.2, 309.1, 309.3, 308.2, 308.5, 307.8, 306.4, 
    306.5, 306.2, 307.5, 309.6, 310.1,
  NaNf, 304.6, 305.1, 310, 309.6, 309.8, 310.6, 310.5, 308.4, 306.9, 307, 
    307.1, 310, 309.5, 309.6, 307.8,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1792, 290.8492, 
    289.7092, 288.8292, 286.1693, 287.2592, 290.8792,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4193, 291.3092, 
    292.0992, 290.6292, 289.2092, 293.0392, 293.1592,
  NaNf, 288.6693, 287.9892, 288.3893, 286.0492, 286.5192, 287.3292, 289.4092, 
    288.8392, 287.5792, 287.4592, 289.3992, 290.6792, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1393, 289.4492, 292.5592, 294.6492, 292.1292, 288.4193, 
    294.1792, 296.4292, 296.1693, 294.5892, 293.3992, 293.8992, NaNf, NaNf,
  NaNf, NaNf, 290.1192, 296.4193, 292.8292, 294.6093, 290.6292, 292.3392, 
    292.6192, 295.1192, 298.0492, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1892, 295.5592, 294.5892, 295.2592, 297.3893, 296.5992, 
    293.0492, 293.8593, 302.8392, NaNf, NaNf, NaNf, 298.5492, NaNf,
  NaNf, 293.2292, 293.5592, 294.9292, 296.7092, 295.0392, 297.6693, 297.1892, 
    296.1292, 297.1093, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6292, 293.7692, 294.5592, 295.5492, 299.1093, 296.6292, 
    296.3792, 299.9392, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.4992, 296.4592, 295.2592, 296.3392, 302.1592, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8492, 
    300.8692, 300.9292, 301.4392, 299.7292,
  NaNf, NaNf, NaNf, NaNf, 298.5492, 296.1892, 300.5192, 301.9892, 301.5992, 
    302.0192, 301.4392, 300.2792, 301.3893, 302.4792, 301.1792, 303.3893,
  NaNf, NaNf, NaNf, NaNf, 300.0692, 301.9492, 300.4392, 301.3792, 302.6592, 
    301.0892, 302.9092, 301.6992, 300.4492, 303.5492, 304.7392, 305.9892,
  NaNf, NaNf, 299.5392, 300.5692, 301.9392, 297.3792, 303.8092, 299.9992, 
    300.6192, 301.3392, 302.6393, 303.6892, 304.4592, 304.6693, 305.6093, 
    306.6093,
  NaNf, 301.1592, 303.8593, 303.1992, 295.6892, 301.8492, 303.0992, 305.7392, 
    303.9992, 305.2892, 305.0092, 305.3992, 305.6192, 305.5992, 306.3992, 
    307.1093,
  NaNf, 298.2992, 297.8893, 303.5892, 302.7492, 307.0592, 307.0692, 306.1992, 
    306.5892, 306.0592, 304.8292, 304.8292, 304.9092, 305.6693, 307.2492, 
    307.4792,
  NaNf, 303.6892, 303.4692, 308.0992, 307.6592, 307.3392, 308.1093, 308.0192, 
    306.6892, 305.7092, 305.6792, 305.7792, 307.6292, 307.2092, 307.1492, 
    305.9792,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.743, 288.613, 
    287.183, 287.373, 284.643, 285.933, 287.873,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.163, 289.543, 
    288.533, 287.063, 287.063, 290.003, 288.953,
  NaNf, 287.813, 287.093, 287.263, 284.563, 285.023, 285.703, 287.773, 
    287.323, 286.443, 286.473, 287.803, 288.503, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.243, 287.523, 289.043, 290.873, 287.673, 286.953, 290.923, 
    292.043, 291.223, 291.933, 289.823, 291.103, NaNf, NaNf,
  NaNf, NaNf, 288.413, 293.543, 288.453, 290.473, 286.933, 289.093, 290.213, 
    292.203, 294.823, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.943, 293.533, 290.673, 291.423, 293.953, 292.483, 289.153, 
    291.083, 301.393, NaNf, NaNf, NaNf, 293.823, NaNf,
  NaNf, 290.643, 290.313, 290.593, 293.243, 291.453, 294.333, 293.813, 
    291.663, 294.293, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.913, 291.913, 291.373, 291.663, 294.113, 292.133, 293.693, 
    296.193, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.363, 292.183, 291.243, 293.873, 299.123, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.343, 
    297.803, 297.893, 298.553, 296.963,
  NaNf, NaNf, NaNf, NaNf, 295.573, 292.413, 297.803, 299.083, 298.373, 
    299.253, 298.063, 297.123, 298.543, 299.623, 298.693, 300.673,
  NaNf, NaNf, NaNf, NaNf, 296.743, 299.973, 297.593, 298.713, 299.873, 
    298.403, 300.213, 299.113, 297.743, 300.773, 301.563, 302.883,
  NaNf, NaNf, 297.133, 298.183, 298.313, 295.413, 301.333, 297.943, 298.383, 
    298.963, 300.033, 300.883, 301.473, 301.703, 302.493, 303.383,
  NaNf, 299.213, 301.713, 300.063, 294.383, 299.743, 300.613, 302.843, 
    301.253, 302.423, 302.143, 302.513, 302.683, 302.703, 303.173, 303.813,
  NaNf, 295.203, 296.343, 301.263, 300.443, 304.093, 304.023, 303.213, 
    304.083, 303.163, 302.293, 302.363, 303.063, 302.993, 303.993, 304.193,
  NaNf, 301.573, 301.003, 305.023, 304.593, 304.153, 304.893, 304.733, 
    304.193, 303.903, 303.823, 303.843, 304.343, 304.013, 303.943, 303.513,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.8925, 292.1925, 
    291.9925, 290.4925, 287.4925, 288.6925, 292.8925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.8925, 292.7925, 
    293.6925, 292.2925, 289.8925, 292.7925, 294.5925,
  NaNf, 289.2925, 288.0925, 287.5925, 283.6925, 283.5925, 286.4925, 289.3925, 
    289.6925, 287.9925, 287.3925, 291.1925, 291.9925, NaNf, NaNf, NaNf,
  NaNf, NaNf, 286.6925, 285.1925, 289.8925, 290.5925, 289.2925, 286.1925, 
    290.2925, 294.0925, 294.3925, 292.5925, 293.4925, 296.2925, NaNf, NaNf,
  NaNf, NaNf, 288.4925, 292.4925, 290.2925, 290.5925, 287.7925, 289.4925, 
    288.2925, 291.5925, 296.2925, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.5925, 292.1925, 292.3925, 292.1925, 293.1925, 291.8925, 
    291.1925, 291.0925, 300.1925, NaNf, NaNf, NaNf, 299.2925, NaNf,
  NaNf, 293.7925, 293.6925, 294.3925, 294.3925, 293.1925, 294.1925, 293.7925, 
    295.3925, 295.4925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.5925, 293.2925, 294.7925, 295.2925, 297.0925, 293.9925, 
    293.6925, 300.0925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 296.0925, 294.6925, 293.8925, 295.0925, 299.1925, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.9925, 
    298.6925, 299.3925, 300.5925, 300.6925,
  NaNf, NaNf, NaNf, NaNf, 294.8925, 295.6925, 297.1925, 299.7925, 298.3925, 
    297.5925, 299.0925, 297.3925, 299.2925, 300.4925, 299.5925, 304.3925,
  NaNf, NaNf, NaNf, NaNf, 296.1925, 297.1925, 297.3925, 297.7925, 298.6925, 
    297.8925, 299.7925, 299.2925, 298.2925, 300.8925, 303.2925, 306.2925,
  NaNf, NaNf, 295.2925, 295.3925, 297.6925, 293.7925, 300.0925, 296.7925, 
    297.1925, 297.4925, 298.6925, 300.9925, 302.3925, 302.6925, 305.2925, 
    307.6925,
  NaNf, 296.5925, 297.4925, 299.0925, 291.5925, 298.3925, 300.5925, 303.1925, 
    300.6925, 302.2925, 303.2925, 304.6925, 305.0925, 304.4925, 306.2925, 
    307.5925,
  NaNf, 295.7925, 293.4925, 299.7925, 298.6925, 305.3925, 304.6925, 303.1925, 
    303.7925, 304.5925, 305.0925, 304.7925, 305.6925, 305.5925, 306.5925, 
    307.4925,
  NaNf, 298.0925, 299.5925, 305.3925, 305.7925, 306.0925, 306.7925, 306.3925, 
    306.1925, 306.2925, 306.2925, 306.7925, 307.3925, 306.4925, 306.8925, 
    306.8925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.9062, 292.4562, 
    291.1963, 289.9662, 287.2362, 288.2863, 292.5562,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.1762, 292.7563, 
    294.8163, 293.2362, 290.4862, 294.3662, 295.3662,
  NaNf, 289.0763, 288.3863, 288.7662, 286.4962, 286.9763, 288.3163, 290.5463, 
    289.9763, 288.4163, 288.2563, 290.6462, 292.1762, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.3763, 289.2362, 293.5463, 295.3163, 293.4062, 289.0262, 
    295.2563, 298.5162, 298.2263, 295.5862, 295.0363, 295.8863, NaNf, NaNf,
  NaNf, NaNf, 290.4362, 296.5463, 293.9362, 295.4362, 291.9163, 293.3563, 
    293.2563, 296.3263, 299.6462, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.4662, 295.6562, 295.5463, 296.0162, 298.1562, 297.3662, 
    294.6462, 294.7762, 303.4262, NaNf, NaNf, NaNf, 300.7062, NaNf,
  NaNf, 294.4562, 294.9163, 296.5562, 297.3062, 295.9763, 298.3362, 298.2563, 
    298.2362, 298.9062, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.1162, 294.4262, 295.9962, 297.2462, 300.8962, 298.1963, 
    298.0463, 302.3763, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.4662, 298.1462, 297.2563, 297.7462, 303.8062, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.7662, 
    302.8362, 303.1063, 303.5862, 302.0162,
  NaNf, NaNf, NaNf, NaNf, 299.1063, 298.1762, 302.0862, 303.9662, 303.0963, 
    303.0963, 303.4562, 302.0862, 303.3763, 304.3863, 302.8563, 305.5262,
  NaNf, NaNf, NaNf, NaNf, 301.0262, 301.8062, 302.0862, 302.8163, 304.0162, 
    302.4763, 304.4362, 303.4763, 302.3062, 305.2762, 307.0162, 308.4662,
  NaNf, NaNf, 299.9262, 300.9662, 303.0162, 298.4862, 304.9262, 301.0862, 
    301.9662, 302.5663, 304.0663, 305.3263, 306.3263, 306.5562, 307.6963, 
    309.2062,
  NaNf, 301.5663, 303.9962, 303.9463, 296.3263, 303.1663, 304.5562, 307.4362, 
    305.5063, 306.8062, 306.6663, 307.2362, 307.5262, 307.5063, 308.6562, 
    309.6462,
  NaNf, 299.7963, 298.9062, 305.1862, 303.9662, 308.9163, 309.0562, 308.0063, 
    308.1862, 307.7162, 306.3763, 306.4362, 306.1462, 307.4662, 309.4763, 
    309.9862,
  NaNf, 304.3163, 304.9763, 309.8163, 309.4862, 309.6063, 310.4262, 310.3163, 
    308.2462, 306.8662, 306.8863, 307.0763, 309.8662, 309.3763, 309.4062, 
    307.7662,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1785, 290.8585, 
    289.7185, 288.8285, 286.1785, 287.2685, 290.8985,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4285, 291.3185, 
    292.1185, 290.6485, 289.2185, 293.0385, 293.1685,
  NaNf, 288.6685, 287.9885, 288.3785, 286.0385, 286.5185, 287.3285, 289.4085, 
    288.8485, 287.5785, 287.4685, 289.4085, 290.6885, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1185, 289.4285, 292.5485, 294.6185, 292.1185, 288.4185, 
    294.1685, 296.4285, 296.1685, 294.5885, 293.4085, 293.9085, NaNf, NaNf,
  NaNf, NaNf, 290.1185, 296.3985, 292.8185, 294.5885, 290.6185, 292.3285, 
    292.6085, 295.1085, 298.0485, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1785, 295.5385, 294.5785, 295.2385, 297.3785, 296.5685, 
    293.0385, 293.8485, 302.8385, NaNf, NaNf, NaNf, 298.5585, NaNf,
  NaNf, 293.2285, 293.5485, 294.9185, 296.6885, 295.0285, 297.6485, 297.1785, 
    296.1285, 297.1085, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.6185, 293.7685, 294.5585, 295.5385, 299.0985, 296.6185, 
    296.3885, 299.9485, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.4885, 296.4485, 295.2585, 296.3385, 302.1585, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8585, 
    300.8785, 300.9385, 301.4585, 299.7385,
  NaNf, NaNf, NaNf, NaNf, 298.5285, 296.1785, 300.5285, 301.9985, 301.5985, 
    302.0085, 301.4485, 300.2785, 301.3985, 302.4885, 301.1885, 303.3985,
  NaNf, NaNf, NaNf, NaNf, 300.0485, 301.9185, 300.4485, 301.3785, 302.6585, 
    301.0885, 302.9085, 301.7085, 300.4585, 303.5585, 304.7485, 306.0085,
  NaNf, NaNf, 299.5285, 300.5485, 301.9185, 297.3785, 303.8085, 299.9985, 
    300.6185, 301.3385, 302.6385, 303.6885, 304.4585, 304.6785, 305.6185, 
    306.6285,
  NaNf, 301.1385, 303.8385, 303.1885, 295.6985, 301.8485, 303.0985, 305.7385, 
    303.9985, 305.2885, 305.0085, 305.4085, 305.6285, 305.6085, 306.4085, 
    307.1185,
  NaNf, 298.2985, 297.8985, 303.5985, 302.7485, 307.0685, 307.0785, 306.2085, 
    306.5985, 306.0585, 304.8285, 304.8285, 304.9085, 305.6785, 307.2585, 
    307.4985,
  NaNf, 303.6785, 303.4685, 308.0985, 307.6685, 307.3485, 308.1185, 308.0285, 
    306.6985, 305.7085, 305.6885, 305.7885, 307.6385, 307.2185, 307.1585, 
    305.9885,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.753, 288.623, 
    287.193, 287.383, 284.653, 285.943, 287.883,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.173, 289.553, 
    288.543, 287.073, 287.073, 290.013, 288.963,
  NaNf, 287.823, 287.093, 287.273, 284.573, 285.033, 285.713, 287.783, 
    287.333, 286.453, 286.483, 287.813, 288.513, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.243, 287.533, 289.053, 290.883, 287.683, 286.963, 290.933, 
    292.053, 291.243, 291.953, 289.843, 291.113, NaNf, NaNf,
  NaNf, NaNf, 288.423, 293.553, 288.463, 290.483, 286.943, 289.113, 290.223, 
    292.213, 294.833, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.953, 293.543, 290.683, 291.433, 293.963, 292.493, 289.163, 
    291.093, 301.393, NaNf, NaNf, NaNf, 293.843, NaNf,
  NaNf, 290.643, 290.323, 290.603, 293.253, 291.463, 294.343, 293.823, 
    291.673, 294.303, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.923, 291.923, 291.383, 291.673, 294.123, 292.143, 293.703, 
    296.203, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.363, 292.193, 291.253, 293.883, 299.143, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.363, 
    297.813, 297.913, 298.563, 296.983,
  NaNf, NaNf, NaNf, NaNf, 295.583, 292.423, 297.813, 299.093, 298.383, 
    299.263, 298.073, 297.143, 298.563, 299.633, 298.703, 300.683,
  NaNf, NaNf, NaNf, NaNf, 296.753, 299.973, 297.613, 298.733, 299.883, 
    298.413, 300.233, 299.133, 297.753, 300.783, 301.573, 302.893,
  NaNf, NaNf, 297.133, 298.193, 298.323, 295.423, 301.343, 297.953, 298.393, 
    298.973, 300.043, 300.903, 301.483, 301.713, 302.513, 303.403,
  NaNf, 299.213, 301.713, 300.073, 294.383, 299.753, 300.623, 302.853, 
    301.263, 302.433, 302.163, 302.533, 302.693, 302.723, 303.183, 303.823,
  NaNf, 295.213, 296.343, 301.273, 300.453, 304.103, 304.033, 303.223, 
    304.093, 303.173, 302.303, 302.373, 303.073, 303.013, 304.003, 304.213,
  NaNf, 301.573, 301.013, 305.033, 304.603, 304.173, 304.913, 304.753, 
    304.203, 303.913, 303.833, 303.853, 304.353, 304.033, 303.963, 303.523,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.2, 292.6, 292, 
    290.7, 287.9, 289, 293.6,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293, 293.8, 296.2, 
    293.5, 290.6, 294.6, 295.7,
  NaNf, 289.8, 289, 288.6, 285.3, 285.1, 287.9, 290.9, 290.8, 288.9, 288.1, 
    291.6, 292.9, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287, 285.9, 292.1, 295.8, 293.4, 287.7, 296.1, 298.8, 298.6, 
    295.7, 296, 297.9, NaNf, NaNf,
  NaNf, NaNf, 288.5, 292.9, 291.8, 293.5, 290.2, 292.3, 291.7, 295.2, 298.5, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 290.1, 294, 294.3, 294.6, 297.2, 296.2, 294.3, 295.6, 306.2, 
    NaNf, NaNf, NaNf, 303.2, NaNf,
  NaNf, 295.9, 295.1, 296.4, 297.1, 295.3, 298.6, 298.2, 298.6, 300, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 298.3, 294.8, 296.6, 298, 301.4, 298.2, 300.1, 306, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 301.2, 299.3, 298.7, 300, 308, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 310.4, 
    306.5, 307.9, 308.6, 306.9,
  NaNf, NaNf, NaNf, NaNf, 300.5, 299.9, 305.8, 308.6, 307.2, 307.4, 307.5, 
    306.1, 307, 308, 307.9, 310.6,
  NaNf, NaNf, NaNf, NaNf, 302.3, 303.6, 305, 306.6, 307, 305.3, 307.8, 307, 
    305.5, 308.3, 311.2, 313.8,
  NaNf, NaNf, 301.3, 301.2, 305.3, 301, 307.7, 304.2, 304.6, 305.3, 307, 
    308.1, 309.4, 309.9, 312, 314.8,
  NaNf, 302, 305, 305.4, 298.6, 306.9, 307.3, 310.3, 308.2, 309.1, 309.3, 
    310.8, 310.9, 310.5, 312.3, 313.4,
  NaNf, 302.1, 301.9, 308.7, 306.6, 312.8, 311.5, 310.3, 311.7, 310.3, 309.3, 
    309.7, 309.7, 311.2, 313.2, 314.2,
  NaNf, 307.1, 307.4, 312.7, 313.5, 312.7, 313.2, 313.4, 310.9, 309.8, 310.1, 
    310.6, 313.3, 313, 313.7, 312.2,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.8, 292.4, 291.2, 
    289.9, 287.2, 288.3, 292.5,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.1, 292.7, 294.7, 
    293.1, 290.4, 294.3, 295.3,
  NaNf, 289.1, 288.4, 288.7, 286.4, 286.9, 288.3, 290.5, 290, 288.4, 288.2, 
    290.6, 292.2, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.3, 289.1, 293.4, 295.1, 293.2, 288.9, 295.1, 298.3, 298, 
    295.4, 294.9, 295.8, NaNf, NaNf,
  NaNf, NaNf, 290.4, 296.3, 293.8, 295.2, 291.8, 293.3, 293.1, 296.1, 299.5, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.4, 295.5, 295.4, 295.9, 298, 297.2, 294.5, 294.6, 303.3, 
    NaNf, NaNf, NaNf, 300.6, NaNf,
  NaNf, 294.4, 294.9, 296.5, 297.2, 295.9, 298.2, 298.1, 298.1, 298.8, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297, 294.4, 295.9, 297.2, 300.7, 298.1, 297.9, 302.2, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.4, 298.1, 297.2, 297.7, 303.7, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.6, 
    302.7, 303, 303.5, 302,
  NaNf, NaNf, NaNf, NaNf, 299, 298.1, 301.9, 303.9, 302.9, 302.9, 303.3, 
    301.9, 303.2, 304.3, 302.8, 305.5,
  NaNf, NaNf, NaNf, NaNf, 300.8, 301.6, 301.9, 302.7, 303.8, 302.3, 304.3, 
    303.3, 302.2, 305.2, 306.9, 308.4,
  NaNf, NaNf, 299.8, 300.8, 302.7, 298.3, 304.8, 300.9, 301.8, 302.4, 303.9, 
    305.2, 306.2, 306.4, 307.6, 309.2,
  NaNf, 301.4, 303.8, 303.7, 296.2, 303, 304.4, 307.3, 305.4, 306.7, 306.6, 
    307.1, 307.4, 307.4, 308.6, 309.6,
  NaNf, 299.7, 298.7, 305, 303.8, 308.8, 308.8, 307.8, 308, 307.6, 306.3, 
    306.4, 306.1, 307.4, 309.4, 309.9,
  NaNf, 304.1, 304.8, 309.7, 309.4, 309.4, 310.2, 310.1, 308.1, 306.8, 306.8, 
    307, 309.7, 309.3, 309.3, 307.7,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1793, 290.8693, 
    289.7193, 288.8393, 286.1793, 287.2693, 290.9193,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4293, 291.3293, 
    292.1193, 290.6593, 289.2193, 293.0392, 293.1893,
  NaNf, 288.6693, 287.9792, 288.3793, 286.0293, 286.5092, 287.3293, 289.4193, 
    288.8593, 287.5893, 287.4693, 289.4193, 290.6992, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.1093, 289.3993, 292.5293, 294.5992, 292.0992, 288.4093, 
    294.1593, 296.4193, 296.1593, 294.5793, 293.3993, 293.9093, NaNf, NaNf,
  NaNf, NaNf, 290.1093, 296.3693, 292.7993, 294.5692, 290.6193, 292.3192, 
    292.5992, 295.1093, 298.0392, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1693, 295.5193, 294.5593, 295.2193, 297.3593, 296.5493, 
    293.0392, 293.8393, 302.8192, NaNf, NaNf, NaNf, 298.5593, NaNf,
  NaNf, 293.2193, 293.5493, 294.8993, 296.6693, 295.0092, 297.6293, 297.1593, 
    296.1193, 297.1093, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.5992, 293.7592, 294.5493, 295.5392, 299.0893, 296.6093, 
    296.3793, 299.9492, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.4693, 296.4393, 295.2592, 296.3393, 302.1593, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8492, 
    300.8793, 300.9393, 301.4593, 299.7493,
  NaNf, NaNf, NaNf, NaNf, 298.5092, 296.1793, 300.5193, 301.9993, 301.5893, 
    301.9893, 301.4492, 300.2693, 301.4093, 302.4993, 301.1893, 303.4093,
  NaNf, NaNf, NaNf, NaNf, 300.0392, 301.8693, 300.4492, 301.3793, 302.6493, 
    301.0793, 302.9093, 301.7093, 300.4593, 303.5593, 304.7592, 306.0193,
  NaNf, NaNf, 299.5092, 300.5293, 301.8993, 297.3793, 303.8093, 299.9993, 
    300.6193, 301.3293, 302.6393, 303.6893, 304.4693, 304.6793, 305.6293, 
    306.6393,
  NaNf, 301.1293, 303.8192, 303.1693, 295.6893, 301.8492, 303.0992, 305.7393, 
    303.9993, 305.2892, 305.0092, 305.4093, 305.6293, 305.6093, 306.4093, 
    307.1293,
  NaNf, 298.2993, 297.8993, 303.5992, 302.7393, 307.0692, 307.0793, 306.2093, 
    306.5992, 306.0593, 304.8393, 304.8393, 304.9193, 305.6793, 307.2693, 
    307.5092,
  NaNf, 303.6593, 303.4693, 308.0992, 307.6693, 307.3593, 308.1193, 308.0293, 
    306.6992, 305.7093, 305.6893, 305.7993, 307.6393, 307.2193, 307.1693, 
    305.9993,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.753, 288.633, 
    287.203, 287.393, 284.663, 285.953, 287.893,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.173, 289.563, 
    288.553, 287.083, 287.083, 290.023, 288.973,
  NaNf, 287.823, 287.103, 287.283, 284.583, 285.033, 285.713, 287.793, 
    287.343, 286.463, 286.483, 287.823, 288.523, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.253, 287.533, 289.063, 290.893, 287.693, 286.973, 290.943, 
    292.063, 291.253, 291.963, 289.853, 291.123, NaNf, NaNf,
  NaNf, NaNf, 288.433, 293.553, 288.473, 290.493, 286.953, 289.123, 290.233, 
    292.223, 294.843, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.953, 293.543, 290.693, 291.443, 293.973, 292.503, 289.173, 
    291.103, 301.393, NaNf, NaNf, NaNf, 293.853, NaNf,
  NaNf, 290.653, 290.323, 290.613, 293.253, 291.473, 294.353, 293.833, 
    291.683, 294.313, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.923, 291.933, 291.393, 291.683, 294.133, 292.153, 293.713, 
    296.213, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.373, 292.203, 291.263, 293.893, 299.153, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.373, 
    297.833, 297.923, 298.583, 296.993,
  NaNf, NaNf, NaNf, NaNf, 295.583, 292.433, 297.823, 299.103, 298.393, 
    299.273, 298.093, 297.153, 298.573, 299.653, 298.713, 300.693,
  NaNf, NaNf, NaNf, NaNf, 296.763, 299.973, 297.623, 298.743, 299.893, 
    298.423, 300.243, 299.143, 297.763, 300.803, 301.583, 302.913,
  NaNf, NaNf, 297.143, 298.203, 298.333, 295.433, 301.353, 297.963, 298.403, 
    298.983, 300.053, 300.913, 301.503, 301.723, 302.523, 303.413,
  NaNf, 299.223, 301.723, 300.083, 294.393, 299.753, 300.633, 302.863, 
    301.273, 302.453, 302.173, 302.543, 302.713, 302.733, 303.203, 303.843,
  NaNf, 295.223, 296.353, 301.283, 300.463, 304.123, 304.043, 303.233, 
    304.113, 303.193, 302.313, 302.383, 303.083, 303.023, 304.023, 304.223,
  NaNf, 301.583, 301.023, 305.043, 304.613, 304.183, 304.923, 304.763, 
    304.213, 303.923, 303.843, 303.863, 304.363, 304.043, 303.973, 303.533,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 294.1925, 293.8925, 
    292.7925, 290.7925, 288.3925, 289.4925, 294.1925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 294.3925, 294.8925, 
    297.6925, 294.9925, 291.7925, 295.9925, 296.4925,
  NaNf, 290.5925, 290.0925, 289.6925, 287.3925, 286.9925, 289.3925, 292.4925, 
    291.9925, 289.7925, 288.9925, 292.4925, 294.0925, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.8925, 286.8925, 294.0925, 298.2925, 296.0925, 289.3925, 
    297.8925, 301.6925, 300.4925, 297.4925, 297.9925, 298.7925, NaNf, NaNf,
  NaNf, NaNf, 288.9925, 295.1925, 293.6925, 297.3925, 292.2925, 295.4925, 
    294.9925, 299.0925, 301.9925, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.3925, 297.0925, 297.1925, 297.8925, 301.2925, 300.1925, 
    297.3925, 298.6925, 305.0925, NaNf, NaNf, NaNf, 304.7925, NaNf,
  NaNf, 298.6925, 296.8925, 299.1925, 300.6925, 298.1925, 302.2925, 301.8925, 
    301.8925, 303.1925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 302.5925, 297.8925, 300.1925, 301.3925, 305.3925, 301.9925, 
    303.0925, 308.2925, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 305.6925, 302.9925, 302.3925, 303.0925, 310.3925, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 313.1925, 
    309.4925, 310.2925, 310.9925, 308.8925,
  NaNf, NaNf, NaNf, NaNf, 303.4925, 303.9925, 309.0925, 311.5925, 309.2925, 
    309.0925, 310.2925, 309.2925, 309.9925, 309.9925, 309.1925, 312.4925,
  NaNf, NaNf, NaNf, NaNf, 306.9925, 306.7925, 309.0925, 309.9925, 310.8925, 
    308.7925, 309.6925, 309.3925, 308.2925, 311.5925, 313.4925, 316.3925,
  NaNf, NaNf, 305.5925, 306.0925, 309.2925, 303.6925, 312.5925, 307.6925, 
    308.3925, 308.8925, 310.5925, 311.4925, 312.6925, 312.9925, 314.5925, 
    316.9925,
  NaNf, 307.8925, 310.9925, 311.0925, 302.3925, 309.9925, 311.2925, 314.3925, 
    311.9925, 313.0925, 312.7925, 313.6925, 313.8925, 313.5925, 314.9925, 
    315.8925,
  NaNf, 307.3925, 306.9925, 313.3925, 307.1925, 317.0925, 315.6925, 314.7925, 
    315.5925, 313.8925, 312.3925, 312.9925, 312.2925, 313.8925, 316.1925, 
    316.7925,
  NaNf, 313.0925, 312.5925, 317.1925, 318.0925, 317.2925, 317.5925, 317.8925, 
    314.4925, 312.4925, 313.2925, 313.6925, 316.1925, 316.0925, 316.5925, 
    314.7925,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.8, 292.4, 291.1, 
    289.9, 287.2, 288.2, 292.5,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.1, 292.7, 294.7, 
    293.1, 290.4, 294.3, 295.2,
  NaNf, 289.1, 288.4, 288.7, 286.4, 286.9, 288.3, 290.5, 289.9, 288.4, 288.2, 
    290.6, 292.2, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.2, 289, 293.4, 295.3, 293.3, 288.9, 295.2, 298.4, 298.1, 
    295.5, 294.9, 295.8, NaNf, NaNf,
  NaNf, NaNf, 290.3, 296.2, 293.8, 295.3, 291.8, 293.3, 293.1, 296.2, 299.5, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.4, 295.6, 295.4, 295.9, 298.1, 297.2, 294.6, 294.8, 303.8, 
    NaNf, NaNf, NaNf, 300.8, NaNf,
  NaNf, 294.5, 294.9, 296.5, 297.3, 295.9, 298.3, 298.2, 298.2, 298.9, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.2, 294.5, 296, 297.2, 300.9, 298.1, 298.1, 302.5, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.6, 298.1, 297.3, 297.8, 304, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.9, 
    302.9, 303.3, 303.8, 302.2,
  NaNf, NaNf, NaNf, NaNf, 299.1, 298.2, 302.2, 304.2, 303.3, 303.4, 303.6, 
    302.2, 303.5, 304.5, 303.1, 305.7,
  NaNf, NaNf, NaNf, NaNf, 301.1, 302.2, 302.2, 303, 304.2, 302.7, 304.5, 
    303.6, 302.4, 305.4, 307.2, 308.6,
  NaNf, NaNf, 300.1, 301, 303.2, 298.7, 305.1, 301.2, 302.1, 302.7, 304.2, 
    305.4, 306.4, 306.7, 307.8, 309.4,
  NaNf, 301.6, 304, 304.1, 296.5, 303.3, 304.7, 307.6, 305.6, 306.8, 306.7, 
    307.4, 307.6, 307.5, 308.7, 309.7,
  NaNf, 299.8, 299.1, 305.3, 304, 309.2, 309.2, 308.1, 308.4, 307.7, 306.4, 
    306.5, 306.2, 307.5, 309.5, 310.1,
  NaNf, 304.5, 305, 309.9, 309.7, 309.8, 310.6, 310.4, 308.3, 306.9, 306.9, 
    307.1, 309.9, 309.5, 309.6, 307.8,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1785, 290.8685, 
    289.7185, 288.8485, 286.1885, 287.2785, 290.9285,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4285, 291.3385, 
    292.1385, 290.6685, 289.2285, 293.0385, 293.1985,
  NaNf, 288.6585, 287.9785, 288.3685, 286.0285, 286.5085, 287.3285, 289.4185, 
    288.8585, 287.5885, 287.4785, 289.4185, 290.6985, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.0885, 289.3785, 292.5185, 294.5685, 292.0885, 288.4085, 
    294.1485, 296.4185, 296.1485, 294.5785, 293.4085, 293.9185, NaNf, NaNf,
  NaNf, NaNf, 290.0985, 296.3285, 292.7785, 294.5485, 290.5985, 292.3085, 
    292.5885, 295.0985, 298.0385, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1585, 295.4985, 294.5485, 295.1985, 297.3285, 296.5185, 
    293.0285, 293.8385, 302.8185, NaNf, NaNf, NaNf, 298.5685, NaNf,
  NaNf, 293.2185, 293.5485, 294.8985, 296.6485, 294.9985, 297.5985, 297.1485, 
    296.1185, 297.1185, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.5885, 293.7485, 294.5385, 295.5285, 299.0785, 296.5985, 
    296.3885, 299.9485, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.4585, 296.4385, 295.2485, 296.3385, 302.1585, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8485, 
    300.8785, 300.9585, 301.4685, 299.7685,
  NaNf, NaNf, NaNf, NaNf, 298.4885, 296.1785, 300.5285, 302.0085, 301.5785, 
    301.9785, 301.4485, 300.2685, 301.4085, 302.5085, 301.1985, 303.4185,
  NaNf, NaNf, NaNf, NaNf, 300.0185, 301.8385, 300.4485, 301.3785, 302.6485, 
    301.0785, 302.9085, 301.7185, 300.4685, 303.5585, 304.7685, 306.0385,
  NaNf, NaNf, 299.4885, 300.5085, 301.8785, 297.3785, 303.7985, 299.9985, 
    300.6285, 301.3285, 302.6385, 303.6885, 304.4685, 304.6885, 305.6285, 
    306.6585,
  NaNf, 301.1185, 303.7985, 303.1485, 295.6885, 301.8485, 303.0985, 305.7385, 
    303.9885, 305.2885, 305.0085, 305.4085, 305.6285, 305.6185, 306.4185, 
    307.1485,
  NaNf, 298.2885, 297.8985, 303.6085, 302.7385, 307.0785, 307.0885, 306.2085, 
    306.5985, 306.0585, 304.8385, 304.8385, 304.9185, 305.6885, 307.2785, 
    307.5185,
  NaNf, 303.6485, 303.4685, 308.0885, 307.6685, 307.3685, 308.1285, 308.0385, 
    306.6985, 305.7185, 305.6885, 305.7985, 307.6485, 307.2285, 307.1785, 
    306.0085,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.763, 288.643, 
    287.213, 287.403, 284.673, 285.963, 287.903,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.183, 289.573, 
    288.563, 287.093, 287.093, 290.033, 288.983,
  NaNf, 287.833, 287.113, 287.293, 284.583, 285.043, 285.723, 287.803, 
    287.353, 286.463, 286.493, 287.833, 288.533, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.263, 287.543, 289.073, 290.913, 287.703, 286.983, 290.953, 
    292.073, 291.263, 291.973, 289.863, 291.133, NaNf, NaNf,
  NaNf, NaNf, 288.433, 293.563, 288.483, 290.503, 286.963, 289.133, 290.243, 
    292.243, 294.853, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.963, 293.553, 290.703, 291.453, 293.983, 292.513, 289.183, 
    291.113, 301.393, NaNf, NaNf, NaNf, 293.863, NaNf,
  NaNf, 290.663, 290.333, 290.623, 293.263, 291.483, 294.363, 293.843, 
    291.693, 294.323, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.933, 291.943, 291.403, 291.693, 294.143, 292.163, 293.723, 
    296.223, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.383, 292.213, 291.273, 293.903, 299.163, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.393, 
    297.843, 297.943, 298.593, 297.003,
  NaNf, NaNf, NaNf, NaNf, 295.593, 292.443, 297.843, 299.113, 298.403, 
    299.283, 298.103, 297.173, 298.583, 299.663, 298.733, 300.703,
  NaNf, NaNf, NaNf, NaNf, 296.763, 299.963, 297.633, 298.753, 299.913, 
    298.443, 300.253, 299.153, 297.783, 300.813, 301.603, 302.923,
  NaNf, NaNf, 297.153, 298.213, 298.343, 295.443, 301.363, 297.973, 298.413, 
    298.993, 300.063, 300.923, 301.513, 301.743, 302.533, 303.423,
  NaNf, 299.233, 301.733, 300.093, 294.403, 299.763, 300.643, 302.873, 
    301.283, 302.463, 302.183, 302.553, 302.723, 302.743, 303.213, 303.853,
  NaNf, 295.233, 296.353, 301.293, 300.473, 304.133, 304.053, 303.253, 
    304.123, 303.203, 302.323, 302.393, 303.093, 303.033, 304.033, 304.233,
  NaNf, 301.583, 301.033, 305.063, 304.623, 304.193, 304.933, 304.783, 
    304.223, 303.933, 303.853, 303.873, 304.383, 304.063, 303.993, 303.553,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.9, 292.6, 291.9, 
    289.9, 287.1, 288.1, 292.8,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.3, 294, 295.8, 
    293.6, 290.2, 294.3, 294.6,
  NaNf, 290.1, 289.5, 289, 286.4, 285.7, 288.1, 290.6, 290.6, 288.7, 287.9, 
    291.8, 292.7, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.9, 286.9, 292.3, 294.4, 293.2, 288.8, 295.2, 298.9, 298.4, 
    295.1, 295.3, 296.4, NaNf, NaNf,
  NaNf, NaNf, 289.2, 293.8, 292, 294.8, 291, 293.5, 292.2, 294.8, 298.2, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1, 295.4, 296.3, 296.9, 298.4, 297, 294.5, 294.4, 301.5, 
    NaNf, NaNf, NaNf, 301.1, NaNf,
  NaNf, 296.9, 295.9, 297.5, 298.4, 296.4, 298.5, 298.2, 298.9, 299.1, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 298.3, 296.8, 298.4, 299.2, 301.9, 298.4, 297.9, 303, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 301.4, 299.5, 298.3, 298.1, 303.1, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.2, 
    303.8, 303.7, 304.6, 303.3,
  NaNf, NaNf, NaNf, NaNf, 298.9, 299.7, 301.8, 304.2, 302.9, 302.3, 303.9, 
    302.8, 303.8, 304.6, 303.3, 307.6,
  NaNf, NaNf, NaNf, NaNf, 301.1, 301.5, 302.3, 302.3, 303.6, 302.4, 304.4, 
    304.1, 303, 307.1, 307.2, 310,
  NaNf, NaNf, 299.6, 300.2, 303.5, 298, 306, 300.9, 302.2, 303, 304.2, 305.8, 
    306.7, 307.1, 308.8, 311,
  NaNf, 302.1, 303.4, 304.8, 296.2, 302.9, 305.2, 307.9, 305.4, 307.3, 307.5, 
    308.1, 309.1, 308.5, 310.1, 310.9,
  NaNf, 301.5, 299.1, 305.8, 301.4, 308.4, 308.7, 308.3, 308.8, 308.9, 308.5, 
    308.8, 308.5, 309.5, 311.4, 311.8,
  NaNf, 304.9, 306.1, 311.1, 310.4, 310.1, 310.6, 311.2, 310.2, 309.6, 309.6, 
    309.9, 311.2, 311.1, 311.4, 310.1,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.8, 292.3, 291.1, 
    289.9, 287.2, 288.2, 292.4,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 293.1, 292.7, 294.7, 
    293.1, 290.4, 294.3, 295.2,
  NaNf, 289.1, 288.4, 288.7, 286.4, 286.9, 288.2, 290.5, 289.9, 288.3, 288.2, 
    290.6, 292.1, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.2, 289, 293.4, 295.3, 293.3, 288.9, 295.2, 298.5, 298.1, 
    295.5, 295, 295.8, NaNf, NaNf,
  NaNf, NaNf, 290.3, 296.2, 293.7, 295.3, 291.7, 293.3, 293.1, 296.2, 299.5, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.4, 295.6, 295.4, 295.9, 298.1, 297.2, 294.6, 294.8, 303.6, 
    NaNf, NaNf, NaNf, 300.8, NaNf,
  NaNf, 294.5, 294.9, 296.5, 297.4, 295.9, 298.4, 298.2, 298.2, 298.9, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 297.4, 294.5, 296, 297.2, 300.9, 298.1, 298.1, 302.5, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 299.7, 298.2, 297.3, 297.8, 304, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 306.9, 
    302.9, 303.3, 303.8, 302.2,
  NaNf, NaNf, NaNf, NaNf, 299.2, 298.2, 302.4, 304.3, 303.4, 303.5, 303.7, 
    302.3, 303.6, 304.6, 303.2, 305.7,
  NaNf, NaNf, NaNf, NaNf, 301.2, 302.3, 302.4, 303.1, 304.3, 302.8, 304.6, 
    303.7, 302.4, 305.4, 307.2, 308.7,
  NaNf, NaNf, 300.2, 301, 303.3, 298.8, 305.2, 301.3, 302.1, 302.8, 304.3, 
    305.5, 306.5, 306.7, 307.9, 309.5,
  NaNf, 301.7, 304.2, 304.3, 296.6, 303.4, 304.7, 307.7, 305.7, 306.9, 306.8, 
    307.4, 307.7, 307.6, 308.8, 309.8,
  NaNf, 300, 299.3, 305.5, 303.9, 309.3, 309.3, 308.1, 308.5, 307.8, 306.4, 
    306.6, 306.2, 307.6, 309.6, 310.1,
  NaNf, 304.7, 305.1, 309.9, 309.7, 309.9, 310.7, 310.5, 308.3, 306.9, 307, 
    307.1, 310, 309.5, 309.6, 307.9,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.1693, 290.8792, 
    289.7292, 288.8492, 286.1892, 287.2892, 290.9492,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 292.4292, 291.3392, 
    292.1393, 290.6792, 289.2392, 293.0392, 293.2092,
  NaNf, 288.6592, 287.9792, 288.3692, 286.0192, 286.4992, 287.3292, 289.4193, 
    288.8692, 287.5892, 287.4692, 289.4292, 290.7092, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.0792, 289.3593, 292.4992, 294.5492, 292.0692, 288.3992, 
    294.1393, 296.4092, 296.1393, 294.5692, 293.4092, 293.9292, NaNf, NaNf,
  NaNf, NaNf, 290.0892, 296.2992, 292.7692, 294.5292, 290.5892, 292.2992, 
    292.5692, 295.0892, 298.0392, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 291.1592, 295.4692, 294.5292, 295.1792, 297.3192, 296.4892, 
    293.0192, 293.8292, 302.8192, NaNf, NaNf, NaNf, 298.5892, NaNf,
  NaNf, 293.2192, 293.5392, 294.8893, 296.6292, 294.9792, 297.5792, 297.1292, 
    296.1093, 297.1192, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 296.5692, 293.7492, 294.5392, 295.5292, 299.0592, 296.5892, 
    296.3893, 299.9592, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 298.4492, 296.4292, 295.2492, 296.3392, 302.1592, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 304.8492, 
    300.8893, 300.9692, 301.4892, 299.7792,
  NaNf, NaNf, NaNf, NaNf, 298.4792, 296.1792, 300.5292, 302.0192, 301.5792, 
    301.9792, 301.4492, 300.2792, 301.4193, 302.5092, 301.2092, 303.4392,
  NaNf, NaNf, NaNf, NaNf, 300.0092, 301.8292, 300.4492, 301.3792, 302.6492, 
    301.0792, 302.9092, 301.7292, 300.4792, 303.5692, 304.7792, 306.0592,
  NaNf, NaNf, 299.4792, 300.4892, 301.8692, 297.3792, 303.7992, 299.9992, 
    300.6292, 301.3292, 302.6393, 303.6992, 304.4692, 304.6892, 305.6393, 
    306.6792,
  NaNf, 301.1093, 303.7792, 303.1393, 295.6892, 301.8593, 303.0992, 305.7392, 
    303.9992, 305.2892, 305.0192, 305.4193, 305.6393, 305.6192, 306.4292, 
    307.1592,
  NaNf, 298.2892, 297.9092, 303.6192, 302.7392, 307.0892, 307.0992, 306.2192, 
    306.6192, 306.0692, 304.8392, 304.8492, 304.9292, 305.6892, 307.2792, 
    307.5292,
  NaNf, 303.6492, 303.4792, 308.0992, 307.6693, 307.3792, 308.1492, 308.0492, 
    306.7092, 305.7192, 305.6992, 305.8092, 307.6592, 307.2392, 307.1892, 
    306.0192,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 290.773, 288.643, 
    287.223, 287.413, 284.683, 285.973, 287.913,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 291.183, 289.583, 
    288.573, 287.103, 287.103, 290.043, 288.993,
  NaNf, 287.833, 287.113, 287.303, 284.593, 285.053, 285.733, 287.813, 
    287.353, 286.473, 286.503, 287.833, 288.543, NaNf, NaNf, NaNf,
  NaNf, NaNf, 287.273, 287.553, 289.083, 290.923, 287.723, 286.993, 290.963, 
    292.083, 291.273, 291.983, 289.873, 291.143, NaNf, NaNf,
  NaNf, NaNf, 288.443, 293.573, 288.493, 290.513, 286.973, 289.143, 290.253, 
    292.253, 294.863, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 289.963, 293.553, 290.713, 291.463, 293.993, 292.523, 289.193, 
    291.123, 301.383, NaNf, NaNf, NaNf, 293.873, NaNf,
  NaNf, 290.663, 290.343, 290.623, 293.273, 291.493, 294.373, 293.853, 
    291.703, 294.333, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, 293.943, 291.943, 291.403, 291.703, 294.153, 292.173, 293.743, 
    296.243, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, 295.393, 292.223, 291.283, 293.913, 299.173, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf,
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 301.403, 
    297.853, 297.963, 298.603, 297.023,
  NaNf, NaNf, NaNf, NaNf, 295.603, 292.453, 297.853, 299.133, 298.423, 
    299.293, 298.123, 297.183, 298.593, 299.673, 298.743, 300.713,
  NaNf, NaNf, NaNf, NaNf, 296.773, 299.963, 297.653, 298.763, 299.923, 
    298.453, 300.263, 299.163, 297.793, 300.823, 301.613, 302.933,
  NaNf, NaNf, 297.153, 298.223, 298.353, 295.453, 301.373, 297.983, 298.423, 
    299.003, 300.073, 300.933, 301.523, 301.753, 302.553, 303.443,
  NaNf, 299.233, 301.733, 300.103, 294.403, 299.773, 300.653, 302.883, 
    301.303, 302.473, 302.193, 302.563, 302.733, 302.753, 303.233, 303.863,
  NaNf, 295.243, 296.363, 301.303, 300.483, 304.143, 304.073, 303.263, 
    304.133, 303.213, 302.343, 302.403, 303.103, 303.053, 304.053, 304.253,
  NaNf, 301.593, 301.043, 305.073, 304.633, 304.213, 304.953, 304.793, 
    304.233, 303.933, 303.863, 303.883, 304.393, 304.073, 304.003, 303.563 ;

 LatLon_181X360-0p50S-180p00E = _ ;
}
