netcdf CF_H.5.1.2 {
  dimensions:
      station = 5;
      pressure = 3;
      time = 4;
      name_strlen = 3;
  variables:
      char station_name(station, name_strlen);
        station_name:cf_role = "timeseries_id";
        station_name:long_name = "station name";

      float temperature(station, time, pressure);
        temperature:standard_name = "air_temperature";
        temperature:coordinates = "lat lon time pressure station_name";
        temperature:units = "K" ;

      double time(time);
        time:standard_name = "time";
        time:long_name = "time of measurement";
        time:units = "hours since 2019-01-01 00:00:00";

      float lon(station);
        lon:standard_name = "longitude" ;
        lon:long_name = "station longitude";
        lon:units = "degrees_east";
        lon:axis = "X" ;

      float lat(station);
        lat:standard_name = "latitude" ;
        lat:long_name = "station latitude";
        lat:units = "degrees_north";
        lat:axis = "Y" ;

      float pressure(pressure);
        pressure:standard_name = "air_pressure";
        pressure:long_name = "pressure";
        pressure:units = "hPa";
        pressure:axis = "Z";

  // global attributes:
  :featureType = "timeSeriesProfile";
  :Conventions = "CF-1.6";

  data:
    station_name = "AAA", "BBB", "CCC", "DDD", "EEE" ;
    time = 0.0, 12.0, 24.0, 48.0 ;
    lon = -150.5, -105.0, -73.3, -3.5, 97.46 ;
    lat = 61.5, 40.0, 42.5, 50.6, 16.85 ;
    pressure = 1000.0, 850.0, 500.0 ;

    temperature = 273.15, 274.0, 275.0,
                  276.0, 277.0, 278.0,
                  278.1, 278.2, 278.3,
                  278.4, 279.0, 279.1,

                  279.2, 276.3, 276.4,
                  280.0, 280.1, 280.2,
                  280.3, 280.4, 281.0,
                  281.1, 281.2, 281.3,

                  281.4, 282.0, 282.1,
                  282.2, 282.3, 282.4,
                  283.0, 283.1, 283.2,
                  283.3, 283.4, 284.0,

                  284.1, 284.2, 284.3,
                  284.4, 285.0, 285.1,
                  285.2, 285.3, 285.4,
                  286.0, 286.1, 286.2,

                  286.4, 287.0, 287.1,
                  287.2, 287.3, 287.4,
                  288.0, 288.1, 288.3,
                  288.4, 289.0, 289.1 ;


}