netcdf CAMPS_StnProfile_PressureLevels {
   dimensions:
     station = 5 ; // 2584 ;
     stn_name_strlen = 4 ;
     time = 2 ;
     pressure_level = 6 ;

   variables:
     double reftime ;
       reftime:units = "hours since 2019-08-14T18:00:00Z" ;
       reftime:standard_name = "forecast_reference_time" ;
       reftime:long_name = "reference time" ;
       reftime:calendar = "proleptic_gregorian" ;
     double time(time) ;
       time:standard_name = "time";
       time:long_name = "time of measurement" ;
       time:units = "hours since 2019-08-14T18:00:00Z" ;
       time:calendar = "proleptic_gregorian" ;
     float lon(station) ;
       lon:standard_name = "longitude";
       lon:long_name = "station longitude";
       lon:units = "degrees_east";
     float lat(station) ;
       lat:standard_name = "latitude";
       lat:long_name = "station latitude" ;
       lat:units = "degrees_north" ;
     char station_name(station, stn_name_strlen) ;
       station_name:standard_name = "platform_id" ;
       station_name:long_name = "ICAO METAR call letters" ;
       station_name:comment = " Only currently archives reports from stations only if the first letter of the ICAO ID is \'K\', \'P\', \'M\', \'C\', or \'T\'. " ;
       station_name:cf_role = "timeseries_id";

     float pressure_level(pressure_level) ;
       pressure_level:standard_name = "air_pressure" ;
       pressure_level:units = "hPa" ;
       pressure_level:positive = "down" ;
       pressure_level:axis = "Z" ;

     float Temp_instant(station, time, pressure_level) ;
         Temp_instant:standard_name = "air_temperature" ;
         Temp_instant:units = "K" ;
         Temp_instant:coordinates = "time lat lon pressure_level station_name" ;

     float DewPt_instant(station, time, pressure_level) ;
         DewPt_instant:standard_name = "dew_point_temperature" ;
         DewPt_instant:units = "K" ;
         DewPt_instant:coordinates = "time lat lon pressure_level station_name" ;

     float RelHum_instant(station, time, pressure_level) ;
         RelHum_instant:standard_name = "relative_humidity" ;
         RelHum_instant:coordinates = "time lat lon pressure_level station_name" ;

   // global attributes
       :featureType = "timeSeriesProfile";
       :Conventions = "CF-1.6";


   data:
       reftime = 0.0 ;
       time = 0.0, 3.0 ;
       pressure_level = 1000., 975., 950., 925., 850., 700 ;

       lat = 45.8667, 44.0198, 37.7667, 30.2167, 42.89 ; //, 41.1008, 61.93, 43.4167, 43.65, 33.4204, 44.75, 49.1833, 45.8833, 65.2833, 39.1625, 19.97, 34.2167, 43.0, 55.15, 21.4167, 21.62, 48.05, 38.286, 66.07, 52.1833, 55.75, 51.8833, 61.8643, 59.05, 38.8983, 57.75, 53.9, 51.1, 53.63, 41.3, 61.3667, 37.0667, 49.2167, 69.73, 42.57, 34.3, 40.7473, 34.2568, 46.45, 38.9949, 34.0998, 41.8678, 34.75, 40.75, 33.63, 27.495, 32.9667, 41.7, 33.6225, 38.8167, 30.3667, 39.4039, 35.82, 42.885, 34.7325, 40.2247, 36.5833, 30.9018, 21.15, 35.21, 27.3953, 33.4667, 35.4881, 35.8333, 34.5975, 28.85, 42.63, 47.5, 31.2667, 40.8731, 45.4968, 39.9, 38.38, 30.7353, 41.3497, 45.6, 52.12, 46.45, 45.82, 61.1333, 49.45, 54.58, 50.7, 30.22, 51.8667, 50.1833, 48.3667, 49.3833, 49.2, 52.85, 39.0667, 42.0625, 45.0, 49.41, 33.8, 44.02, 41.6, 31.8575, 39.53, 45.65, 32.5117, 47.4542, 48.8844, 41.8756, 41.45, 33.14, 41.1958, 37.2667, 18.4333, 28.1003, 34.8833, 31.4213, 44.68, 36.0167, 48.7837, 41.6333, 35.8497, 41.33, 41.9333, 35.4726, 30.6118, 35.65, 43.72, 36.8553, 35.3333, 36.0833, 41.5261, 34.9, 32.6566, 34.9, 40.7833, 40.1667, 40.8264, 38.5018, 36.3667, 43.1167, 41.2102, 37.3167, 24.55, 33.3, 35.1667, 31.05, 36.77, 48.3008, 34.6018, 39.8333, 37.9333, 39.7, 61.75, 69.6667, 58.42, 44.43, 61.25, 48.9357, 49.1667, 58.4167, 69.62, 44.05, 42.4333, 59.933, 64.9333, 43.0833, 31.7794, 37.2863, 34.67, 32.8683, 53.5833, 61.1, 33.8333, 49.2167, 44.2233, 55.35, 70.32, 64.32, 55.58, 28.7333, 53.6667, 40.67, 30.9167, 35.44, 41.25, 40.3147, 43.6833, 38.9306, 31.5833, 35.14, 32.2153, 32.4667, 34.7229, 31.3275, 38.01, 42.1667, 44.9403, 40.8192, 35.3333, 47.45, 31.8692, 34.65, 47.84, 34.81, 46.1189, 29.5667, 50.1833, 46.54, 48.45, 39.45, 46.15, 33.7172, 36.7667, 47.85, 34.2997, 34.6833, 42.7317, 49.0333, 36.6167, 36.3, 39.2167, 30.3431, 38.0667, 42.4222, 48.5144, 37.1333, 41.1833, 47.25, 41.74, 34.47, 33.94, 31.4667, 35.8579, 60.1667, 46.99, 46.5333, 31.1522, 47.7167, 33.9667, 47.7912, 48.47, 29.3333, 38.6, 66.8175, 42.7275, 31.554, 52.7719, 40.4833, 29.48, 44.5833, 36.35, 44.0167, 39.1333, 34.7167, 38.1833, 41.45, 30.4833, 34.7893, 34.65, 35.2435, 34.1283, 59.5167, 40.4561, 56.65, 42.1, 20.7856, 45.95, 21.4333, 49.9167, 52.9333, 32.5667, 52.1833, 46.1167, 42.2, 56.33, 45.1961, 40.8, 33.9167, 40.4833, 44.45, 41.5097, 37.6333, 40.6306, 38.3566, 37.0318, 45.01, 29.2667, 33.4939, 36.6646, 39.3667, 33.65, 42.9667, 37.3, 34.75, 46.9167, 43.1333, 44.8833, 44.9331, 41.7, 29.9833, 42.2497, 56.9667, 30.4667, 29.5333, 40.92, 45.1667, 33.0375, 39.5, 36.7367, 42.993, 42.7955, 40.9333, 47.5, 40.0833, 32.8875, 45.55, 27.2, 38.27, 49.0833, 46.68, 46.21, 60.77, 45.7, 32.6167, 44.7873, 39.2833, 41.7333, 36.9062, 54.9167, 51.1667, 45.72, 41.02, 41.68, 41.81, 34.2291, 37.8, 40.0972, 36.2, 41.1167, 44.9167, 37.3667, 44.3667, 27.195, 33.27, 32.8525, 30.2906, 35.0333, 33.65, 35.1575, 38.3667, 32.9, 42.2333, 27.9667, 30.4, 37.4167, 46.8333, 33.2, 32.53, 41.89, 33.11, 45.43, 40.1998, 38.5315, 48.3114, 32.6986, 29.9469, 36.45, 30.4, 31.5333, 47.2167, 36.03, 41.8, 33.2856, 30.3925, 30.2436, 35.1351, 48.7754, 32.5645, 42.4, 45.7833, 43.3333, 49.0333, 60.7167, 54.4667, 43.0333, 66.15, 47.7, 53.8833, 50.1167, 50.0167, 20.9, 53.5667, 52.1667, 49.6167, 39.7, 58.3667, 34.65, 35.6697, 33.5977, 41.828, 31.8457, 56.32, 29.6342, 59.727, 32.8292, 34.6905, 33.6333, 66.5667, 32.9733, 47.2899, 49.1, 35.0206, 35.2333, 40.5167, 38.9667, 37.0911, 43.7764, 40.7289, 32.6091, 42.8, 34.4333, 51.9333, 43.65, 40.6069, 41.78, 46.6186, 70.4673, 46.1442, 39.6014, 44.55, 45.43, 55.83, 44.2833, 43.1655, 28.6, 33.9667, 32.7419, 44.4803, 27.7678, 37.2833, 37.6142, 45.78, 34.9157, 39.8333, 34.2, 48.8, 33.6186, 36.5333, 40.18, 37.2978, 38.3106, 41.4833, 49.0167, 41.3302, 38.55, 39.2833, 44.4167, 65.5667, 50.33, 53.4333, 46.67, 25.6419, 28.29, 31.429, 46.8156, 29.805, 45.4182, 31.6659, 42.4667, 34.0225, 46.0229, 38.0972, 44.08, 36.3989, 39.22, 33.5871, 40.62, 45.1167, 44.5833, 31.0425, 34.056, 32.646, 30.5979, 29.9667, 43.1083, 38.95, 34.85, 37.6167, 36.61, 44.35, 36.28, 47.95, 34.6452, 18.57, 39.645, 39.0158, 26.5333, 43.9167, 48.7833, 32.51, 38.8667, 36.29, 37.9333, 33.1783, 44.3333, 40.05, 42.9, 28.0002, 34.7667, 33.95, 45.5511, 40.9502, 35.3167, 48.1833, 26.2456, 42.7586, 44.3667, 44.4042, 45.97, 40.7953, 35.95, 34.6333, 65.2833, 27.8118, 47.16, 48.7667, 45.3, 45.17, 51.67, 47.28, 40.5694, 68.32, 50.7, 50.3833, 46.0106, 38.7167, 49.3, 66.976, 58.1853, 63.7326, 59.75, 66.0, 46.7, 43.98, 59.324, 30.47, 40.0333, 44.0511, 50.7, 65.6226, 41.5667, 33.3667, 27.65, 28.8673, 53.3333, 39.2748, 37.2333, 49.7, 38.85, 40.35, 42.85, 38.9806, 33.8285, 55.2833, 50.25, 56.3667, 34.7333, 32.9549, 42.05, 30.1945, 39.7833, 44.9272, 41.8833, 45.4167, 40.9, 32.6151, 35.9403, 43.67, 37.0639, 46.25, 42.5694, 44.8333, 37.4064, 38.6833, 18.05, 12.2, 12.15, 12.5, 41.5333, 17.48, 45.28, 40.7667, 33.8167, 33.0167, 37.2392, 41.7333, 31.3667, 46.2206, 37.5167, 36.9377, 27.95, 46.39, 42.3667, 32.5792, 37.9833, 39.1333, 42.5429, 55.7, 30.7833, 42.0746, 43.5667, 36.5728, 32.85, 30.0333, 46.4119, 39.0005, 34.8536, 29.1833, 38.9767, 44.0219, 47.4667, 45.07, 39.9461, 39.9, 43.2781, 43.55, 27.655, 43.6833, 48.6, 49.4167, 53.3167, 58.75, 50.2833, 56.8667, 48.65, 46.2833, 49.4667, 58.8333, 54.8167, 51.1167, 46.3667, 41.2261, 29.2111, 30.5271, 37.6333, 30.6833, 48.2553, 43.62, 53.7667, 45.57, 41.34, 38.7815, 38.5393, 41.6667, 46.4267, 31.5367, 52.3597, 29.9, 42.4833, 47.104, 53.6333, 39.25, 45.5644, 38.6065, 38.4333, 46.0167, 49.75, 45.7805, 48.7667, 50.2667, 46.22, 43.42, 35.9373, 47.8, 36.3792, 49.5, 49.49, 29.35, 40.4812, 30.52, 43.95, 40.45, 47.08, 45.8986, 44.5333, 43.43, 51.18, 37.6004, 29.12, 17.1167, 42.03, 30.3833, 43.29, 70.77, 18.5, 17.9333, 46.1667, 34.3833, 31.1062, 45.3, 39.05, 29.3419, 36.3175, 34.4167, 44.5, 36.8933, 40.1522, 36.6886, 35.1333, 29.3667, 35.4333, 32.3372, 44.3333, 36.6167, 41.3333, 30.8317, 37.15, 34.2256, 37.1584, 38.1433, 45.2333, 35.75, 44.61, 39.9, 41.6167, 34.4031, 34.2667, 45.1833, 42.6133, 37.5587, 28.5767, 48.95, 33.0678, 29.6167, 38.9548, 48.55, 26.1775, 47.2833, 44.9833, 55.3, 43.0, 45.25, 53.25, 50.2167, 50.6833, 50.6, 55.3, 41.59, 45.6194, 45.8833, 41.5725, 47.6458, 37.3333, 35.6128, 58.6836, 62.1883, 65.6979, 59.6333, 59.2439, 39.64, 37.7, 44.5691, 38.91, 48.2667, 68.63, 49.8333, 49.3667, 33.6167, 30.8717, 34.2836, 41.2406, 33.6325, 42.8372, 34.4333, 33.95, 36.0233, 40.8667, 46.768, 37.6667, 39.75, 44.32, 31.8833, 29.95, 38.51, 45.2333, 32.3344, 42.43, 49.7667, 40.7333, 35.9728, 39.0495, 34.3105, 33.902, 37.0637, 31.2336, 37.0833, 30.2, 34.17, 40.65, 66.62, 40.9792, 42.05, 34.72, 47.4167, 31.1106, 35.0222, 36.1167, 40.1994, 41.98, 27.5333, 33.2578, 43.5833, 36.4333, 43.18, 29.91, 39.0167, 67.5667, 55.15, 51.38, 45.4691, 33.18, 44.2491, 34.98, 41.45, 31.4208, 42.68, 38.72, 48.1, 42.2413, 46.9667, 37.65, 43.7747, 41.7833, 39.15, 40.5, 38.55, 41.3167, 42.9333, 35.0667, 40.72, 38.8833, 32.3667, 35.8167, 40.0307, 46.3478, 41.6256, 33.5, 35.25, 48.3904, 41.3072, 35.65, 32.4674, 43.5333, 51.45, 47.9167, 48.9285, 53.8667, 35.4606, 37.4667, 48.7531, 50.3667, 38.7842, 44.15, 32.35, 34.8913, 29.4448, 39.1683, 41.0667, 33.9667, 36.3, 48.4047, 51.7667, 43.63, 44.1167, 31.9513, 41.15, 53.0833, 51.1333, 69.15, 54.09, 64.05, 42.2333, 48.02, 49.12, 48.83, 62.95, 42.1, 66.8667, 56.0075, 35.5333, 27.6927, 46.72, 31.48, 50.27, 48.0667, 58.0961, 47.4833, 64.5119, 60.533, 47.05, 38.7606, 38.1, 46.3833, 44.7366, 46.55, 41.7833, 41.4, 33.6494, 42.3512, 37.8667, 39.0083, 45.15, 42.7167, 30.7833, 40.1167, 40.9, 42.05, 39.65, 32.1951, 38.1417, 43.6212, 41.0254, 47.4394, 30.65, 47.3806, 30.22, 45.94, 33.8578, 44.7833, 44.3667, 48.3518, 45.5481, 41.8333, 36.75, 41.65, 41.28, 50.31, 39.0854, 46.58, 48.17, 37.3333, 26.5842, 31.4767, 43.6333, 28.82, 38.9146, 44.05, 40.15, 38.0333, 32.2167, 32.1667, 43.78, 29.7167, 39.2811, 32.2597, 38.7074, 44.8888, 39.6083, 32.5, 42.1667, 43.9667, 39.1333, 19.75, 35.86, 38.5167, 32.85, 35.6167, 32.7333, 38.15, 29.5333, 46.35, 32.1333, 38.7167, 38.0304, 32.4558, 34.6722, 22.0228, 53.0267, 34.4736, 49.7906, 41.3, 38.25, 48.4614, 45.0667, 48.4167, 25.8167, 32.6989, 40.2333, 46.2667, 34.2667, 43.5167, 42.11, 39.3667, 56.02, 40.63, 54.8475, 55.32, 63.6833, 27.0716, 70.2, 61.72, 62.07, 57.15, 59.4467, 66.27, 57.0667, 68.3, 61.1, 52.1167, 29.47, 37.13, 60.48, 52.7167, 68.1336, 49.5167, 32.921, 41.6042, 32.6833, 43.2333, 47.95, 43.3381, 47.5047, 27.7783, 43.5333, 33.9094, 47.4, 53.3167, 43.45, 69.35, 34.7333, 38.05, 41.275, 55.5333, 54.0197, 40.4818, 66.9167, 37.6308, 45.7596, 38.2638, 34.8486, 35.1806, 40.6, 46.82, 49.1333, 48.42, 34.98, 50.1167, 53.03, 29.6167, 38.9557, 66.9833, 33.9167, 48.6167, 52.4333, 45.35, 54.17, 61.58, 45.95, 51.57, 40.8, 33.6317, 36.8207, 35.8953, 34.1833, 45.8667, 26.0667, 29.5061, 35.1333, 43.77, 39.4667, 43.08, 45.7, 47.5928, 36.422, 35.0, 38.9457, 41.9167, 36.2925, 52.2333, 50.95, 54.7667, 54.3, 48.4167, 54.13, 69.6, 53.92, 43.9833, 50.95, 33.45, 50.2333, 38.8333, 30.68, 33.45, 36.3298, 36.75, 47.4833, 44.05, 35.36, 35.0, 38.3392, 33.6667, 41.3839, 41.1, 44.17, 36.6667, 29.8253, 51.48, 34.18, 46.9112, 34.71, 59.45, 62.65, 55.0333, 42.0667, 42.6894, 36.7801, 41.7333, 61.1697, 61.5833, 34.1681, 64.55, 40.2167, 36.6951, 43.22, 33.3013, 39.4274, 40.85, 44.6833, 43.43, 39.4166, 41.1881, 39.6154, 41.27, 45.57, 32.7692, 33.5695, 33.8977, 49.9, 44.63, 45.6983, 39.2119, 37.7, 36.88, 33.2398, 37.77, 68.12, 38.1333, 49.6642, 36.3167, 61.7749, 32.3833, 36.1737, 64.7272, 42.23, 43.9833, 49.63, 45.07, 33.9667, 47.3228, 43.9667, 34.1203, 30.1314, 42.15, 39.2281, 39.07, 43.52, 45.25, 28.4667, 46.8333, 29.8448, 29.3667, 18.4667, 40.2797, 34.5167, 19.47, 45.07, 56.55, 50.03, 45.7, 46.3, 56.65, 44.6, 49.18, 42.45, 27.2628, 31.7357, 43.03, 43.65, 44.35, 52.19, 48.0167, 46.28, 49.2, 36.5321, 49.9, 47.05, 57.5804, 49.15, 44.75, 57.53, 45.68, 49.57, 46.42, 62.12, 35.5083, 40.65, 35.8494, 44.5447, 45.7066, 35.6352, 38.5339, 30.5155, 36.9333, 26.9185, 56.8167, 43.9667, 33.3, 37.7833, 35.4167, 28.65, 40.1961, 47.2667, 34.9027, 41.7833, 43.8317, 34.86, 40.29, 44.016, 56.58, 32.3833, 45.1, 42.59, 46.5667, 42.9167, 40.7, 46.4503, 53.05, 45.506, 41.6833, 35.0833, 38.05, 46.7439, 50.7083, 46.0486, 60.37, 61.2167, 39.734, 62.0954, 43.1702, 55.1311, 38.2833, 39.6167, 63.8833, 59.4333, 33.912, 62.9561, 41.03, 33.31, 34.3833, 34.5071, 38.9914, 51.4667, 43.87, 43.07, 34.9, 33.535, 33.2544, 39.1, 39.47, 44.8922, 72.0, 36.6667, 43.7333, 49.0236, 47.35, 34.4758, 29.65, 48.3833, 38.0894, 50.7, 49.7833, 35.9499, 44.8667, 47.3978, 49.08, 49.25, 32.6833, 46.43, 31.0559, 43.9333, 33.97, 40.85, 38.66, 36.7, 42.55, 38.95, 47.78, 31.25, 30.1167, 43.5667, 39.8167, 42.2419, 46.84, 37.6, 48.48, 30.2896, 42.5, 41.93, 26.3785, 44.2507, 37.22, 31.307, 40.5703, 37.7022, 32.6453, 41.92, 39.08, 29.5622, 37.5211, 43.98, 35.2, 30.5857, 36.9814, 36.0, 41.0375, 34.2667, 40.9, 35.23, 31.0847, 60.5, 31.25, 61.7833, 55.2208, 61.8453, 32.7561, 43.7792, 38.85, 35.57, 44.99, 31.58, 29.17, 36.9, 35.6, 35.6667, 31.9168, 39.1167, 50.05, 42.95, 43.1667, 33.1855, 44.2167, 42.4708, 33.6833, 38.48, 39.1, 28.2167, 32.8167, 70.22, 33.98, 44.8833, 40.2183, 31.6159, 41.42, 35.0, 44.3156, 34.7914, 35.8667, 35.05, 32.3333, 45.5, 40.3833, 39.1923, 39.9194, 41.02, 34.5454, 44.2667, 44.7531, 30.3567, 36.4042, 32.4442, 47.1333, 31.8333, 47.3081, 34.3, 42.6167, 52.1736, 42.15, 23.1333, 36.9875, 48.31, 61.1167, 46.677, 44.36, 54.2333, 36.3616, 69.03, 27.7667, 33.1333, 32.0311, 38.3667, 47.9167, 49.85, 49.2, 51.4667, 38.2489, 48.4333, 33.8167, 47.57, 30.3333, 42.9667, 42.2333, 55.62, 40.0833, 40.45, 48.9406, 53.55, 55.2, 41.02, 50.55, 47.0, 49.62, 58.7, 45.7667, 50.55, 45.9667, 51.1833, 69.28, 22.15, 40.6839, 49.83, 45.12, 46.84, 53.33, 44.8167, 50.2, 21.35, 44.4833, 46.18, 34.6, 43.9833, 36.93, 35.2891, 31.42, 36.0425, 42.2667, 42.75, 33.7833, 38.8, 38.65, 26.2, 18.0167, 42.6, 27.7411, 31.6072, 32.8333, 38.8833, 42.55, 37.45, 46.1, 32.9147, 43.2348, 44.99, 61.42, 41.35, 36.37, 71.2842, 42.5667, 45.3728, 32.2126, 35.8893, 43.28, 45.1403, 60.7833, 70.1333, 55.2, 39.45, 65.99, 64.0, 37.4495, 37.7, 40.2394, 36.03, 70.3443, 68.8833, 61.18, 37.18, 31.6167, 42.6667, 61.5363, 29.72, 33.2167, 43.5794, 44.0435, 49.9667, 42.1667, 47.0338, 47.8167, 34.65, 30.7506, 19.78, 31.8111, 52.2333, 53.3167, 39.2833, 42.1075, 28.5464, 31.1793, 68.35, 27.835, 42.2667, 56.95, 45.32, 41.9833, 42.5667, 36.9, 30.0692, 48.02, 42.98, 41.4364, 33.3667, 34.6217, 46.4167, 29.248, 27.727, 44.58, 48.7081, 45.67, 56.2333, 53.2167, 58.45, 44.2333, 54.3, 35.1, 58.7667, 37.05, 33.65, 41.1333, 40.2833, 29.1153, 34.98, 33.5931, 34.6, 30.0719, 37.81, 38.7167, 48.2994, 32.0365, 33.9781, 43.0333, 47.9872, 70.17, 35.6558, 33.65, 35.935, 36.63, 44.1333, 41.07, 40.45, 35.2667, 38.9467, 42.6, 39.3333, 39.4833, 24.7262, 38.5, 44.5, 69.4333, 51.15, 48.6, 48.75, 52.35, 34.2667, 53.55, 53.7, 32.6992, 54.28, 36.2, 52.0667, 33.9, 43.05, 46.0093, 44.3931, 37.5, 39.53, 32.7469, 41.2744, 40.8167, 26.1833, 44.6333, 33.7794, 42.3667, 45.65, 37.65, 42.4536, 38.69, 47.6333, 35.0199, 29.5189, 48.85, 30.3564, 43.5667, 33.527, 48.5333, 30.0481, 44.51, 39.5856, 36.77, 46.7, 46.8667, 49.8167, 25.4833, 34.65, 45.6833, 37.95, 36.25, 34.7073, 36.6869, 63.6167, 33.95, 39.95, 40.5, 47.95, 35.2322, 40.9167, 51.2667, 43.8789, 32.3239, 19.7167, 38.7833, 41.4, 24.5757, 42.6431, 41.02, 35.95, 36.2667, 35.35, 35.35, 31.3822, 27.5072, 32.5167, 45.3723, 48.1333, 42.5519, 49.5, 49.89, 32.85, 49.7, 45.37, 49.1167, 41.54, 50.15, 48.27, 52.45, 33.4044, 53.3, 41.0467, 34.5667, 41.3164, 36.0833, 32.552, 33.9333, 40.4167, 38.0667, 42.7833, 20.78, 27.9889, 35.8798, 22.9833, 40.7667, 33.8667, 45.9861, 33.1753, 45.88, 46.9258, 43.7424, 46.7997, 35.2333, 31.5397, 47.2833, 33.995, 30.73, 40.2044, 43.32, 37.0542, 38.7, 41.9906, 34.0136, 45.1167, 61.6, 45.31, 52.2203, 44.5167, 42.7818, 44.9975, 36.2, 28.01, 41.37, 43.65, 32.19, 34.8167, 32.1167, 43.05, 40.4333, 36.68, 70.6392, 42.4667, 67.57, 43.9844, 42.1333, 44.45, 49.3333, 33.0953, 56.4667, 35.72, 44.9167, 40.0833, 61.5717, 34.9915, 42.2667, 38.35, 53.9667, 46.8, 44.9667, 46.1167, 49.6333, 49.7833, 21.4776, 43.8333, 60.1167, 52.7667, 51.2667, 55.1833, 48.3667, 18.3333, 50.4333, 49.7167, 17.7, 37.65, 53.0333, 46.1667, 32.3, 45.43, 41.5092, 33.9167, 36.6541, 39.77, 44.6252, 32.1417, 18.25, 39.5936, 41.75, 39.65, 42.2, 27.913, 26.4419, 44.65, 46.31, 29.9767, 41.2667, 42.0833, 39.1167, 35.48, 43.25, 41.0522, 45.03, 47.63, 26.6833, 44.59, 43.02, 33.8833, 30.3527, 45.6833, 45.5958, 48.5167, 39.3833, 50.2667, 34.2729, 40.1833, 53.62, 36.3712, 53.15, 36.66, 49.07, 46.6, 49.65, 37.45, 32.3538, 31.15, 42.9167, 38.5667, 36.77, 47.71, 35.0333, 48.3694, 37.3333, 40.43, 35.58, 33.1598, 35.1944, 40.2833, 41.7833, 28.6167, 45.6333, 37.751, 46.4794, 38.5383, 45.69, 34.5, 45.15, 33.5906, 31.6839, 43.3497, 37.3592, 43.4393, 42.5833, 32.7009, 34.5186, 37.8596, 50.22, 46.4, 68.7833, 40.7833, 25.9, 40.9479, 45.82, 29.7333, 45.4071, 41.0619, 49.126, 38.7667, 36.35, 34.8578, 42.938, 32.4773, 30.4167, 32.2833, 36.2661, 42.78, 26.2333, 32.8978, 42.595, 45.8258, 39.55, 53.9667, 34.9167, 44.7295, 50.1833, 32.95, 48.7167, 67.73, 55.1163, 61.5408, 45.1177, 25.9, 44.0946, 61.1333, 41.1667, 52.185, 40.0378, 45.62, 41.7092, 35.42, 48.5167, 21.3167, 50.9667, 62.82, 19.9, 39.5803, 36.3333, 30.75, 34.681, 39.7852, 36.0211, 30.7044, 28.2086, 37.9, 37.1667, 33.4667, 32.8167, 42.6167, 33.7833, 31.3183, 60.2, 40.7504, 61.5242, 35.6377, 50.1441, 68.3167, 43.6421, 36.45, 32.6333, 40.0536, 32.0167, 36.4333, 35.76, 35.2167, 25.05, 41.1167, 41.4, 37.7, 36.2117, 44.97, 38.3167, 44.5333, 29.3833, 52.8167, 51.7833, 50.58, 49.4878, 38.1333, 34.4, 50.63, 48.0689, 44.7167, 45.92, 42.25, 35.02, 41.6, 28.0833, 47.75, 35.135, 44.0667, 43.1667, 40.85, 43.6629, 41.69, 49.8344, 35.05, 37.95, 41.07, 44.2667, 42.57, 41.6258, 43.4, 39.8233, 32.6639, 38.8042, 45.75, 31.3833, 43.1143, 36.4129, 33.3117, 41.9167, 46.9, 40.47, 38.05, 34.3093, 38.8167, 28.4533, 38.8167, 45.3167, 33.5294, 43.2, 31.8411, 27.962, 43.9228, 46.9728, 28.2333, 47.7667, 44.5167, 54.4167, 32.4333, 57.5, 30.1692, 46.9, 44.76, 33.7167, 34.7583, 39.35, 33.4167, 28.6539, 30.7167, 41.6167, 58.18, 43.3, 35.0, 44.66, 49.7, 46.35, 43.7667, 44.87, 42.75, 47.83, 54.98, 53.5, 44.66, 41.3833, 50.65, 34.0253, 34.7129, 45.4622, 41.6833, 43.6768, 27.9011, 37.0833, 29.7239, 38.2236, 41.5333, 31.3558, 40.0681, 40.1375, 46.4833, 53.75, 38.38, 41.0, 38.215, 40.16, 44.4755, 37.75, 42.78, 41.1992, 32.5652, 27.9167, 41.4914, 41.5167, 43.1167, 44.28, 41.45, 40.7081, 41.1409, 42.25, 40.2964, 36.2167, 39.1333, 38.3333, 34.81, 47.6333, 40.435, 59.45, 34.2, 49.3372, 33.0634, 42.69, 49.458, 36.03, 40.3331, 58.4167, 66.8881, 50.1289, 46.72, 62.15, 64.55, 63.7833, 42.9333, 64.7333, 50.1014, 49.5263, 41.5, 34.2803, 36.1667, 32.3167, 34.2686, 30.8857, 30.5, 47.7966, 41.1667, 40.3013, 31.85, 43.6, 41.1833, 45.8, 34.5467, 37.3667, 31.3975, 43.92, 32.7822, 42.7461, 44.2667, 47.2, 36.46, 46.7667, 30.4167, 43.1167, 41.6, 36.02, 42.2167, 33.4639, 35.7, 30.9715, 41.12, 46.3036, 40.0228, 63.8833, 42.8667, 44.8, 42.2186, 45.3167, 20.9631, 45.4333, 46.6333, 21.3167, 30.8367, 34.1812, 43.5813, 32.6933, 31.95, 36.98, 41.5631, 36.28, 40.3287, 39.4283, 30.3583, 50.28, 31.0833, 39.6667, 28.9542, 39.531, 44.71, 45.65, 49.25, 37.75, 45.4167, 34.2962, 32.5667, 30.3919, 42.4833, 47.07, 35.66, 68.75, 31.2694, 49.32, 37.5, 45.5, 45.61, 46.35, 38.3154, 27.3496, 45.2667, 54.72, 51.67, 43.8333, 56.55, 45.05, 49.2667, 56.08, 37.1681, 58.3833, 53.6833, 52.82, 50.8167, 50.45, 54.6833, 39.3167, 36.4833, 33.6319, 32.7136, 36.685, 18.5, 34.3155, 49.9058, 45.9658, 51.2, 49.25, 47.5667, 48.6511, 53.03, 34.45, 44.7667, 26.9688, 41.0167, 51.1003, 44.63, 26.15, 41.3461, 39.5639, 68.8, 38.2167, 45.0667, 39.42, 30.5333, 40.78, 44.4667, 63.0186, 61.2667, 41.4148, 41.3667, 67.1, 34.2333, 64.83, 64.8167, 37.0364, 45.9647, 42.3, 18.45, 35.25, 37.0, 28.43, 35.2133, 35.5383, 44.62, 34.3522, 30.5833, 48.1167, 37.82, 41.4, 47.5333, 41.9619, 43.15, 30.6333, 35.4167, 48.15, 41.8, 41.8667, 65.1667, 60.7331, 65.2404, 39.4947, 59.05, 53.8889, 62.3, 44.78, 62.9, 60.79, 55.8, 19.7388, 53.8333, 43.9333, 64.2167, 43.6333, 44.1167, 48.5667, 30.0667, 49.9167, 45.5333, 48.726, 48.2167, 51.4167, 40.1217, 43.2111, 46.5333, 49.1333, 46.154, 40.85, 48.3333, 47.4228, 42.8167, 44.27, 29.229, 36.68, 40.65, 32.9, 32.4167, 42.0458, 41.9167, 45.45, 35.54, 47.6667, 35.05, 37.35, 28.7833, 43.3939, 37.6167, 52.8167, 32.6333, 37.1858, 37.3, 35.6667, 28.5167, 66.2422, 45.55, 33.4331, 56.2333, 46.1731, 44.55, 39.7667, 40.6153, 38.75, 38.5, 44.9333, 31.92, 40.9467, 44.45, 33.5667, 30.9667, 44.2, 39.9406, 41.6167, 41.1389, 34.2667, 47.3833, 49.75, 49.4833, 51.67, 56.37, 49.35, 31.6058, 43.7667, 40.6239, 44.4167, 49.0333, 42.25, 35.93, 50.63, 41.7667, 44.23, 38.3981, 38.2578, 43.2333, 34.35, 33.2333, 35.5448, 38.85, 45.8167, 45.55, 18.27, 40.5167, 44.2667, 33.2333, 47.15, 33.6017, 28.0667, 63.4901, 40.1003, 51.1833, 42.0983, 57.9167, 51.4167, 40.0102, 44.8833, 45.3833, 30.3842, 28.634, 42.9167, 26.1597, 45.1589, 31.4667, 40.6667, 41.9833, 41.94, 44.3814, 40.4915, 45.1, 42.2167, 41.9598, 62.23, 39.3614, 48.5614, 47.8, 37.5136, 38.53, 48.25, 48.3, 30.4967, 68.47, 49.5667, 50.45, 45.5167, 64.7764, 61.25, 45.8333, 60.5667, 62.77, 35.6855, 58.65, 64.65, 67.8167, 40.1637, 30.2358, 48.5572, 37.0906, 34.6, 44.8601, 29.6222, 41.25, 32.1108, 58.9902, 34.045, 35.43, 47.97, 42.4072, 34.0132, 37.2333, 35.3878, 39.8466, 39.8306, 29.2543, 44.0735, 29.97, 39.8333, 42.7, 31.395, 34.2139, 41.7, 45.23, 43.4588, 40.0333, 40.0, 26.0014, 39.05, 40.8217, 35.3055, 30.7836, 38.5863, 37.9, 49.32, 47.1656, 45.24, 36.4372, 30.07, 40.1333, 29.123, 46.2441, 64.78, 39.1833, 36.9667, 31.7936, 35.5977, 31.3167, 43.5, 44.8437, 27.1816, 42.4, 30.5, 38.2667, 33.93, 46.69, 38.65, 31.023, 36.0, 39.7, 32.719, 44.8428, 39.979, 41.9333, 36.7451, 41.5167, 27.2067, 35.9167, 43.4667, 28.4667, 37.7833, 37.0833, 40.52, 44.3, 42.22, 35.2833, 45.31, 28.9731, 37.7355, 44.12, 44.38, 42.1908, 28.96, 42.5417, 21.9833, 47.249, 45.4667, 68.9333, 43.39, 48.2, 35.38, 57.25, 32.48, 35.4, 33.2194, 43.1544, 35.67, 40.5282, 39.15, 38.6667, 31.1819, 37.2848, 45.87, 27.85, 39.3167, 40.2167, 29.714, 37.7416, 28.4333, 32.7, 36.6106, 39.7333, 35.1667, 29.6833, 48.5667, 32.0833, 31.7803, 35.0167, 36.1333, 32.6753, 36.5872, 52.1, 45.22, 44.4333, 34.6988, 40.7333, 61.7603, 32.3667, 35.78, 44.3833, 33.4333, 17.3, 40.4719, 37.1322, 37.7214, 34.9856, 39.8833, 42.9111, 46.07, 54.25, 50.2333, 52.93, 49.08, 53.578, 50.22, 54.15, 50.9, 37.974, 49.3333, 53.1833, 47.3, 60.23, 69.5667, 48.42, 51.3, 49.73, 51.43, 49.0333, 51.0767, 48.4267, 47.4111, 49.68, 50.47, 42.4667, 50.0, 50.23, 43.9752, 20.98, 40.0167, 38.0511, 49.05, 65.22, 31.15, 48.7527, 42.87, 61.25, 27.9156, 32.8344, 54.32, 28.0833, 49.4, 41.7667, 48.88, 51.0833, 45.9, 32.4122, 43.9889, 28.3692, 38.1833, 50.19, 41.2647, 49.63, 46.2833, 41.05, 39.8333, 30.03, 36.1333, 47.97, 36.0167, 33.35, 47.3258, 42.5833, 35.7333, 48.1167, 37.5779, 48.4708, 35.9475, 40.7667, 36.75, 41.7286, 33.6903, 29.3332, 43.9868, 51.0333, 60.1167, 45.8255, 34.2472, 47.0833, 44.4833, 40.9667, 31.0667, 42.8833, 48.3767 ;
       lon = -66.5333, -92.4831, -99.9667, -81.8833, -73.25 ; //, -92.4444, -147.17, -124.25, -95.5833, -112.6862, -81.1, -123.1833, -82.5667, -126.8, -89.6746, -75.85, -118.4833, -82.3, -105.2667, -77.85, -81.55, -77.7833, -76.4118, -162.77, -113.9, -120.1833, -176.65, -162.0261, -158.5167, -119.9947, -152.5167, -166.5333, -100.05, -111.68, -93.12, -139.05, -88.7667, -57.4, -163.02, -84.81, -97.0167, -122.9223, -111.3393, -95.21, -79.1459, -93.0661, -84.0794, -118.7333, -95.42, -91.75, -80.3683, -96.8333, -94.92, -111.9083, -76.8667, -104.0167, -77.975, -81.61, -90.2317, -76.6569, -83.3516, -121.85, -83.8811, -157.1, -91.74, -82.5542, -105.5333, -97.8236, -90.65, -117.383, -96.9167, -83.98, -94.9333, -85.7167, -81.8867, -91.0005, -105.1167, -121.96, -101.203, -71.7989, -103.55, -101.23, -61.97, -73.43, -100.9, -108.9833, -130.7, -120.45, -96.37, -63.2833, -96.0667, -89.1167, -126.55, -113.28, -111.87, -95.6333, -104.1528, -75.63, -82.44, -118.3333, -92.83, -83.8, -86.0108, -89.33, -68.6833, -92.0314, -115.6697, -99.6208, -71.0211, -90.5167, -83.24, -96.1122, -104.3333, -66.0, -80.6356, -95.7833, -97.797, -84.73, -89.4, -97.632, -91.55, -97.4156, -72.045, -72.6833, -98.0053, -81.4612, -109.07, -85.5, -84.8561, -77.9667, -79.95, -85.7867, -120.45, -114.606, -82.2167, -73.9667, -103.2167, -115.7875, -77.3053, -94.1, -77.6667, -81.2516, -79.9667, -81.75, -104.5333, -79.0167, -93.1833, -90.32, -102.4064, -78.5793, -86.3, -75.4667, -77.7167, -121.2333, -121.6667, -130.0, -65.2, -123.75, -57.9104, -105.9667, -130.0, -140.2, -103.0667, -73.3, -164.031, -161.15, -70.8167, -95.7061, -107.056, -120.47, -117.1425, -116.45, -94.07, -116.5, -102.9667, -76.5994, -131.7, -149.58, -158.73, -133.08, -96.25, -113.4667, -91.33, -102.9167, -94.8, -76.9167, -78.8308, -93.3667, -90.4325, -110.3333, -106.8, -98.1777, -93.8167, -80.8546, -92.5486, -77.97, -120.4, -73.0975, -76.8661, -94.3667, -122.3, -95.2172, -98.4, -90.36, -96.67, -67.7939, -90.6667, -61.8, -90.92, -123.3, -87.3, -123.8833, -79.857, -119.7167, -96.62, -90.5123, -86.6833, -95.556, -119.4333, -87.4114, -77.17, -106.8667, -89.8219, -97.8667, -87.8678, -68.4684, -76.6167, -78.9, -123.15, -83.66, -97.96, -96.39, -109.6, -102.0131, -132.75, -94.2, -61.0833, -81.3908, -104.1833, -80.4833, -99.9317, -67.43, -98.4833, -92.1667, -161.0223, -114.4531, -81.8825, -108.2556, -88.9333, -93.63, -71.1833, -94.22, -117.0167, -86.6167, -120.5667, -85.7333, -87.0, -86.5167, -81.1958, -86.94, -97.4708, -84.8472, -139.6667, -106.7403, -111.2167, -83.16, -156.9514, -77.3167, -157.7667, -97.2333, -66.8667, -116.9833, -122.05, -122.9, -72.5333, -103.28, -123.1322, -74.4167, -80.8, -85.6833, -95.8167, -72.8278, -118.85, -93.9008, -93.6842, -85.9537, -84.7, -94.8667, -90.9811, -88.3728, -101.7, -97.2, -79.3333, -108.6333, -87.6167, -114.0833, -89.3333, -93.2167, -74.8492, -74.8, -90.25, -111.3416, -133.95, -87.2, -98.2833, -88.63, -92.5333, -116.9158, -119.7833, -97.1019, -84.1389, -109.8071, -90.4333, -122.2167, -75.0167, -112.72, -93.6, -92.2, -77.45, -61.7, -71.95, -70.79, -137.58, -65.15, -116.4667, -88.56, -80.2333, -72.65, -94.0128, -109.9667, -96.6333, -73.38, -74.73, -93.02, -85.44, -86.2558, -116.7833, -92.5433, -81.65, -111.9667, -97.15, -120.5667, -84.6833, -90.027, -111.82, -104.4675, -97.6958, -85.2, -84.4333, -114.5594, -82.55, -80.0333, -83.3333, -82.5333, -86.47, -122.05, -95.8833, -97.2, -93.75, -89.08, -98.5553, -91.76, -75.1482, -121.7865, -114.2551, -97.0465, -100.1739, -103.15, -89.0667, -81.5333, -93.5167, -76.57, -107.2, -117.4565, -97.5621, -98.9094, -90.2344, -123.1283, -82.9853, -90.7, -111.15, -72.5167, -122.3667, -135.0667, -128.5833, -81.15, -65.72, -79.85, -122.6833, -91.9, -110.7167, -156.4333, -113.5167, -106.6833, -115.7833, -87.67, -134.5833, -112.4333, -120.6283, -83.139, -94.1598, -86.6107, -158.36, -104.3615, -157.259, -115.6717, -77.03, -95.45, -145.2667, -97.3181, -101.581, -123.3, -80.0771, -120.6333, -106.8667, -104.8167, -95.5664, -87.8497, -73.4133, -82.3699, -72.0, -119.8333, -131.0167, -94.4167, -95.8657, -80.7, -93.3097, -157.4357, -115.5964, -116.0056, -110.4167, -73.93, -108.43, -66.3333, -95.2028, -91.2, -98.4833, -95.4964, -103.783, -82.6261, -102.6139, -116.2642, -122.84, -81.9565, -89.6667, -119.2, -122.5333, -114.7142, -115.5667, -74.13, -81.2036, -75.1239, -73.1333, -122.7667, -86.6648, -89.85, -120.7, -72.0167, -167.9167, -105.56, -91.7667, -60.4, -80.4347, -81.44, -83.4885, -74.0939, -95.8979, -123.8144, -98.1486, -98.6833, -106.9031, -92.8952, -106.1686, -91.7, -76.0161, -104.63, -80.2087, -83.06, -87.6333, -124.05, -86.3116, -117.6012, -93.2981, -84.5574, -95.35, -78.9381, -77.45, -82.35, -97.2667, -94.74, -105.5333, -94.31, -97.4, -106.8337, -68.37, -77.468, -87.6497, -81.75, -92.5, -123.05, -92.59, -98.8167, -95.48, -100.7167, -86.7817, -89.0198, -107.88, -72.2667, -82.1642, -114.6167, -117.45, -122.4089, -95.9179, -77.6333, -103.6333, -80.1114, -87.8178, -89.8333, -118.9625, -86.17, -73.1003, -112.15, -118.0833, -126.75, -97.0888, -67.83, -71.7167, -73.35, -73.68, -105.4, -70.63, -102.2727, -100.08, -96.57, -102.5833, -102.6497, -77.5167, -115.1, -160.4365, -157.3856, -148.9106, -154.9167, -153.7, -68.05, -96.32, -155.9018, -88.53, -74.3536, -101.6011, -120.45, -168.0949, -81.4833, -81.9667, -81.3333, -82.5713, -104.01, -103.6659, -89.5833, -86.95, -99.2667, -79.9333, -73.95, -76.9223, -79.1222, -77.7667, -63.6, -94.7, -92.2333, -111.7668, -94.78, -97.6699, -121.85, -89.6242, -91.7, -64.35, -97.98, -85.434, -89.8308, -92.93, -89.2232, -84.4667, -77.7144, -93.45, -77.5248, -104.7667, -63.1167, -68.9667, -68.2833, -70.0167, -93.65, -62.98, -118.0, -73.9, -118.15, -85.0667, -76.7158, -89.6833, -100.5, -100.2456, -122.25, -76.2893, -81.7833, -94.8, -71.0333, -96.7189, -122.05, -75.4667, -83.1779, -119.23, -83.2833, -124.2901, -116.2167, -79.3353, -96.85, -90.0333, -86.6508, -80.2737, -116.7858, -81.05, -76.33, -82.7931, -87.8667, -64.49, -81.8931, -84.2, -70.9222, -80.2167, -80.4142, -79.6333, -68.2, -82.4667, -60.4167, -94.0667, -107.6833, -101.0667, -123.4333, -63.1333, -119.6, -122.6, -127.1833, -114.0167, -79.4167, -92.4939, -99.7433, -98.3588, -120.95, -88.25, -101.2733, -84.74, -125.9833, -95.97, -84.43, -106.2198, -76.0304, -70.2833, -105.8825, -84.1939, -108.8347, -97.87, -76.4667, -122.287, -77.7, -102.28, -84.7928, -87.7267, -113.0167, -91.45, -84.1667, -96.5435, -64.4833, -117.8167, -72.65, -88.13, -77.5465, -69.55, -97.7911, -98.0333, -117.3, -99.1667, -107.2177, -90.42, -78.1667, -99.33, -64.0, -94.8739, -69.6667, -83.86, -112.5, -81.5593, -91.87, -61.7833, -82.9, -84.3667, -79.91, -117.8, -77.9167, -76.7833, -60.05, -103.3167, -98.1959, -85.27, -84.6667, -98.8509, -119.6294, -103.0833, -123.2833, -121.4103, -97.5869, -78.0542, -78.9333, -100.9167, -82.55, -90.2264, -93.3167, -116.0167, -75.7333, -93.3399, -107.75, -99.2836, -95.7784, -122.556, -63.05, -81.3833, -63.42, -83.13, -90.5833, -80.1192, -83.8333, -89.7, -89.59, -82.5674, -94.9767, -95.33, -96.0653, -95.1667, -121.0817, -109.7667, -97.9731, -68.3167, -64.9167, -123.1333, -82.3167, -122.77, -131.8167, -66.2667, -127.3667, -120.5167, -114.7833, -95.34, -121.1714, -82.5667, -86.7345, -101.4394, -95.5167, -100.9961, -156.6539, -159.7749, -156.3514, -151.5, -135.5094, -90.78, -113.1, -72.018, -121.35, -92.4833, -95.85, -92.75, -121.4833, -92.7667, -96.6222, -80.5649, -96.5946, -83.8496, -103.0978, -100.2833, -83.3167, -78.3303, -74.2833, -100.8944, -95.4833, -82.6667, -94.5, -81.5667, -94.0167, -89.09, -81.6333, -104.2519, -93.87, -77.8, -114.0333, -115.1344, -105.5128, -84.4238, -87.3142, -81.7983, -94.75, -76.35, -92.0, -97.12, -73.7833, -160.0, -124.1058, -93.85, -84.87, -68.3167, -93.1533, -76.4625, -86.6833, -87.5956, -95.38, -99.4667, -81.3883, -118.95, -99.5333, -79.4, -96.95, -74.9167, -139.8333, -105.27, -110.35, -89.8057, -96.59, -95.6073, -89.79, -97.35, -110.8458, -91.97, -88.18, -105.5833, -78.3714, -122.9, -97.4167, -98.0386, -111.85, -96.6667, -122.3, -121.3, -122.3167, -71.4333, -118.15, -95.03, -79.85, -95.4, -83.9833, -86.2514, -104.2575, -73.8819, -90.0833, -93.1, -100.0243, -85.0644, -80.5167, -100.4666, -72.95, -116.3333, -122.2833, -103.2973, -94.6667, -77.9649, -122.1167, -98.3937, -114.4167, -93.8029, -103.1, -91.0333, -79.7596, -90.2611, -77.166, -86.1833, -86.0833, -99.7667, -97.3709, -104.2, -116.63, -123.2167, -85.1289, -104.8167, -114.4333, -106.5833, -140.15, -114.45, -139.15, -83.5333, -65.33, -110.47, -72.55, -141.9333, -87.9, -162.6333, -161.1604, -97.6333, -97.2912, -94.38, -97.32, -64.23, -96.1833, -135.4097, -122.7667, -165.4356, -165.114, -109.4667, -87.5989, -92.55, -117.0167, -85.57, -93.68, -124.2333, -95.05, -81.685, -86.2556, -80.4, -95.2117, -89.13, -71.1167, -86.5167, -85.6167, -117.8, -102.8, -106.9167, -81.8696, -76.4292, -96.2158, -80.4134, -65.5978, -86.52, -92.8322, -93.15, -89.26, -98.4904, -89.6667, -71.55, -122.6559, -122.9544, -90.3333, -108.2333, -70.5167, -91.67, -110.09, -76.7594, -72.73, -122.17, -79.2, -81.8625, -82.8603, -72.3167, -81.81, -82.0986, -70.2833, -122.25, -84.6, -80.7, -110.8833, -82.99, -98.05, -76.61, -107.72, -93.1759, -72.2292, -77.0077, -93.6667, -72.7167, -90.7333, -121.4333, -70.55, -98.42, -121.5, -109.6333, -106.0833, -117.1667, -89.7, -98.4667, -87.4, -81.2, -77.1833, -120.4146, -96.9122, -82.8814, -159.7851, -122.5064, -85.7214, -94.3778, -95.9, -78.05, -119.5192, -93.35, -101.35, -80.2833, -94.9486, -85.3833, -119.1167, -116.85, -112.0667, -92.92, -75.0667, -87.68, -79.1, -163.4103, -160.52, -170.5, -82.4403, -148.4667, -157.15, -163.3, -170.2167, -151.7044, -166.05, -135.35, -133.4833, -155.5667, -124.1333, -92.37, -80.68, -151.03, 174.1, -151.7433, -113.9833, -80.6406, -88.0847, -96.8667, -123.3667, -97.1833, -73.6106, -111.1873, -97.6903, -84.0833, -94.8594, -92.5, -113.5833, -65.47, -124.0667, -118.2167, -87.5333, -111.0322, -102.35, -109.1383, -111.4288, -151.5167, -84.3323, -64.2414, -78.8964, -111.7885, -103.6008, -98.4333, -60.66, -112.05, -64.32, -78.36, -127.9333, -112.82, -83.1, -94.3713, -136.2167, -118.3333, -112.3833, -114.9167, -60.98, -131.67, -64.65, -94.35, -107.92, -99.76, -85.1523, -76.0333, -100.4036, -79.7167, -95.3833, -80.15, -95.4769, -111.6667, -88.4864, -76.1667, -94.27, -90.4, -95.7235, -105.2899, -77.98, -104.5699, -88.25, -92.5851, -87.8833, -107.15, -112.0167, -130.6, -123.3167, -108.53, -130.9, -106.07, -80.75, -127.64, -94.0, -121.5833, -94.9, -97.68, -88.5833, -77.6352, -104.5, -111.3667, -75.7333, -96.94, -78.8833, -75.5042, -117.8833, -72.5059, -102.9833, -114.93, -121.6, -90.035, -107.05, -91.9342, -96.8147, -97.22, -157.328, -160.18, -131.5667, -70.2167, -90.4444, -76.4488, -71.4333, -150.0261, -159.5333, -101.7173, -149.0833, -111.7167, -76.1355, -95.83, -117.3552, -101.0466, -77.85, -111.1167, -88.69, -118.701, -103.6774, -78.7609, -95.77, -93.27, -97.4415, -86.0512, -117.6024, -98.2667, -93.23, -110.4408, -82.2293, -121.8167, -91.91, -119.4582, -90.43, -145.57, -91.7667, -93.7328, -119.4, -161.3194, -86.3667, -94.1191, -155.4699, -91.17, -64.6667, -114.48, -66.47, -117.6333, -71.1483, -86.4, -119.121, -93.3761, -79.25, -106.3161, -88.53, -89.77, -112.55, -80.55, -92.1833, -82.0475, -100.7833, -69.67, -83.1148, -83.9833, -70.7, -77.87, -115.2667, -110.72, -92.95, -63.58, -111.2167, -63.52, -98.08, -81.88, -80.8498, -93.0991, -102.52, -94.98, -78.3, -127.47, -64.5, -76.0, -122.68, -93.2005, -109.47, -91.75, -157.572, -88.35, -63.66, -111.57, -96.99, -57.89, -64.77, -136.18, -108.7925, -86.15, -77.8967, -95.0806, -94.9334, -77.3853, -106.933, -96.7041, -111.45, -81.9939, -132.95, -69.7167, -111.6667, -89.25, -97.3833, -89.8, -76.7731, -122.5833, -76.881, -87.75, -111.8061, -86.56, -88.14, -97.0859, -169.67, -94.7167, -90.3, -117.87, -120.5333, -97.3833, -74.1667, -62.5758, -93.33, -91.9811, -70.9667, -77.05, -97.28, -117.1136, -121.2814, -71.25, -166.27, -149.8333, -77.43, -163.6821, -88.725, -131.5781, -104.5167, -110.75, -152.2833, -146.3333, -84.9406, -155.6058, -93.37, -84.77, -89.55, -81.9472, -76.4833, -109.1667, -79.37, -92.62, -117.8667, -112.3832, -97.5806, -84.4333, -106.15, -91.8678, -125.27, -87.5, -103.6167, -95.5983, -70.03, -93.1042, -95.2833, -123.9167, -88.1231, -119.2833, -123.1667, -96.7731, -91.4833, -120.2014, -66.73, -65.33, -103.2, -63.85, -82.7741, -60.0167, -80.99, -72.6333, -88.45, -76.9, -94.1833, -95.6667, -93.65, -82.4, -93.2167, -71.4333, -82.9333, -96.9814, -96.66, -83.3167, -99.2364, -87.6718, -79.28, -88.71, -80.1077, -90.8553, -80.42, -95.4038, -75.4883, -112.1544, -81.5964, -84.59, -77.57, -91.5256, -76.7644, -94.55, -81.15, -100.6486, -77.0011, -94.1667, -81.4669, -110.0, -97.62, -79.4, -83.8031, -145.5, -81.4667, -166.0333, -162.7278, -165.5713, -91.8806, -71.7536, -77.0333, -77.05, -96.18, -94.72, -82.22, -81.35, -88.9167, -95.3667, -98.6003, -94.6, -112.13, -87.9, -86.2333, -80.0362, -93.9167, -93.27, -78.9333, -106.32, -121.5667, -89.6167, -117.15, -150.98, -83.67, -116.1, -76.8556, -91.2972, -88.42, -99.05, -69.7972, -79.3681, -78.7833, -90.0, -88.75, -118.4, -75.9667, -119.7326, -76.8769, -95.27, -94.2027, -121.15, -95.5558, -95.4139, -90.6479, -97.8167, -104.8, -104.8, -119.5147, -103.8, -89.0333, -106.7189, -121.7333, -81.2833, -82.53, -71.13, -122.85, -122.9827, -64.2961, -125.7667, -78.5292, -107.82, -97.5, -117.2833, -96.3989, -81.6, -74.6167, -64.45, -98.9, -90.2, -86.9536, -123.4333, -78.7167, -71.23, -81.5167, -83.7333, -85.55, -118.29, -95.5833, -105.0167, -97.9028, -114.1, -119.4, -89.38, -111.85, -65.45, -113.82, -98.5, -62.6833, -103.65, -81.4833, -115.5667, -119.22, -100.98, -92.901, -64.3, -74.29, -71.2, -104.0, -62.3333, -104.7, -157.9333, -79.55, -72.92, -120.07, -70.95, -121.78, -95.0939, -87.05, -95.9894, -84.4667, -73.8, -118.05, -97.65, -88.9667, -80.1833, -66.5667, -95.23, -98.0247, -110.4281, -106.0, -90.05, -92.4, -105.8667, -118.2833, -85.9628, -93.6241, -85.2, -149.52, -89.15, -92.46, -156.7781, -110.1, -72.7739, -101.5216, -101.0301, -91.73, -79.4028, -161.8, -143.6333, -132.83, -74.5667, -161.12, -145.7333, -94.7311, -98.75, -75.5567, -119.07, -150.9447, -166.1333, -149.97, -77.52, -97.2167, -83.4167, -160.3413, -91.33, -92.8139, -90.8965, -89.304, -119.3833, -76.9, -120.5313, -91.8333, -99.2667, -92.6886, -155.55, -106.3758, -87.8833, -110.0667, -114.85, -77.9844, -81.3358, -99.3239, -166.8, -96.013, -71.8667, -158.6167, -95.65, -87.9, -72.2833, -76.2, -93.8036, -92.87, -96.07, -99.6422, -110.75, -79.7344, -92.8, -88.441, -96.191, -92.48, -122.9103, -61.38, -117.4333, -105.6833, -78.1167, -78.3667, -130.45, -97.97, -111.1167, -100.9667, -101.8167, -100.6833, -79.4, -95.4631, -81.06, -95.0633, -79.07, -83.5736, -88.55, -93.55, -116.56, -102.101, -83.9624, -88.2333, -66.3375, -124.68, -105.1381, -88.45, -79.0658, -80.02, -87.6667, -71.92, -109.5167, -113.95, -92.6827, -82.8333, -76.4167, -88.2833, -81.0514, -107.8833, -80.2167, -133.0167, -121.5, -86.3, -91.6167, -97.03, -88.7667, -64.1, -57.0333, -117.2153, -112.97, -95.9, -111.45, -117.25, -108.45, -83.7439, -74.2028, -77.3333, -107.72, -96.5303, -85.84, -82.5167, -98.2333, -90.1833, -82.8158, -122.8667, -84.52, -75.77, -91.9476, -75.3625, -117.5333, -80.6203, -95.2417, -95.7, -95.008, -96.7333, -112.2953, -58.55, -102.2131, -108.07, -85.8, -98.67, -92.5, -68.0167, -74.53, -80.3833, -86.7667, -74.0333, -79.8167, -115.0333, -77.4452, -77.4828, -135.8667, -81.1167, -91.2, -107.5333, -124.55, -75.6225, -81.4333, -80.65, -91.2528, -84.9826, -155.0667, -104.716, -92.9459, -81.6888, -77.0494, -94.37, -85.0811, -76.1833, -89.8667, -99.2, -103.5106, -97.8097, -84.9333, -94.7466, -69.7167, -71.7558, -112.12, -97.13, -106.1, -112.7833, -71.82, -117.7333, -87.53, -60.05, -70.12, -113.75, -118.4133, -132.7667, -78.4117, -98.4167, -105.6722, -115.1667, -88.5555, -118.4, -86.9333, -102.6833, -84.6, -76.32, -82.0186, -106.2694, -82.4, -111.9667, -117.9667, -95.992, -97.8283, -93.27, -98.6692, -111.0978, -102.7997, -101.7, -82.5075, -121.3333, -80.3613, -98.23, -84.5319, -84.69, -84.6149, -121.6, -93.6189, -118.4556, -113.8833, -149.0833, -92.69, -174.2064, -114.2167, -71.5148, -92.8557, -94.4833, -82.35, -91.15, -70.3167, -82.37, -77.6167, -110.9333, -115.8667, -76.5667, -82.03, -159.9948, -71.2833, -162.98, -88.557, -86.4333, -83.4, -123.1833, -94.9614, -132.3833, -96.82, -123.0, -83.0667, -149.5403, -117.8631, -82.9667, -98.87, -101.1, -71.4, -79.3, -64.6833, -112.8, -94.3667, -158.0443, -66.0833, -128.8167, -108.25, -102.4667, -118.8833, -89.3167, -64.9667, -104.6667, -124.9, -64.8, -122.1167, -122.5167, -60.05, -86.4, -84.91, -74.265, -84.5167, -83.2178, -90.24, -86.2008, -94.8517, -65.6333, -84.2264, -72.1833, -79.9167, -89.1, -97.2115, -98.1294, -73.4667, -85.46, -99.0857, -80.6667, -80.1833, -108.5333, -81.16, -79.2167, -93.6897, -102.02, -65.75, -80.1167, -63.55, -91.12, -84.3, -87.3167, -118.85, -122.6092, -123.0167, -99.8333, -107.7333, -78.715, -80.65, -112.03, -82.1734, -115.12, -76.32, -107.58, -112.0, -109.52, -106.8, -97.4338, -97.7167, -106.4667, -90.15, -80.82, -59.31, -79.5, -89.3272, -121.8167, -104.6333, -79.1, -95.6211, -83.8647, -74.8167, -122.4667, -80.7, -89.45, -82.6367, -84.3572, -106.0486, -85.57, -82.7167, -93.2167, -85.8475, -83.2709, -76.3847, -121.9242, -85.9949, -99.9833, -80.0029, -109.3786, -76.8941, -121.58, -94.1333, -81.25, -91.1167, -97.4333, -87.1826, -92.37, -85.0167, -83.8129, -73.7044, -123.0024, -109.75, -97.9167, -102.3264, -85.0606, -80.7231, -86.6833, -106.9167, -93.1558, -96.2, -97.6667, -79.7829, -87.9381, -119.2611, -97.65, -97.8333, -92.15, -96.266, -61.8167, -84.27, -94.6, -164.55, -162.2662, -165.6009, -95.1304, -80.2833, -121.2002, -146.25, -73.1333, -128.1567, -105.2274, -122.65, -92.7349, -80.15, -72.2667, -157.9167, -118.1833, -92.12, -75.1333, -79.3394, -119.95, -95.58, -90.3467, -104.5431, -102.5478, -87.023, -100.0188, -85.9667, -94.5, -82.0333, -97.35, -123.3667, -84.5167, -85.4439, -154.3, -106.2715, -166.1468, -91.1764, -123.1106, -133.5167, -80.4116, -105.6667, -108.1667, -106.3689, -81.1333, -81.4167, -80.96, -83.4167, -77.4667, -95.9, -70.6167, -77.4333, -115.1958, -95.72, -88.8667, -72.6167, -98.5833, -111.1, -114.6833, -126.93, -123.2994, -78.45, -96.15, -96.98, -69.5556, -66.8, -66.6, -81.9, -94.62, -109.0667, -97.05, -90.35, -118.4392, -69.1167, -79.9333, -74.05, -84.2613, -93.5658, -124.4981, -106.6, -107.9, -87.83, -88.5167, -84.42, -80.2122, -94.75, -93.5792, -97.0958, -76.069, -87.05, -92.3, -89.5315, -100.7516, -79.3196, -70.7333, -71.5, -91.43, -103.5167, -81.6407, -92.2167, -99.2169, -104.7167, -75.6667, -82.5164, -71.5, -99.4036, -93.6708, -78.8833, -123.9303, -80.6, -116.8167, -109.0167, -110.2833, -99.85, -134.5833, -96.98, -95.0667, -94.08, -96.6667, -82.3764, -81.4333, -112.3833, -96.6811, -87.0167, -87.4167, -103.7, -79.8, -105.6667, -63.61, -103.8, -63.1667, -99.3167, -94.38, -93.77, -92.68, -85.43, -130.6333, -63.58, -79.8667, -99.93, -118.2881, -79.957, -69.5953, -70.0, -92.1797, -98.0517, -84.0833, -98.6946, -85.6583, -71.2833, -85.7512, -118.5692, -75.265, -84.51, -73.67, -88.41, -85.2, -83.5874, -89.33, -93.0163, -97.22, -105.37, -74.6261, -97.3081, -82.6833, -120.5644, -88.1833, -76.1167, -85.42, -96.52, -84.0214, -104.8691, -89.58, -78.32, -81.0833, -123.2, -96.2, -82.7029, -117.65, -75.3817, -135.3167, -118.3667, -124.3939, -80.2793, -88.3, -123.7152, -79.47, -75.1222, -135.7333, -157.1624, -122.9547, -92.04, -145.45, -163.03, -171.75, -78.7333, -156.9333, -122.9356, -123.4963, -74.1, -87.6004, -97.0833, -90.0833, -86.8583, -94.0349, -81.7, -103.2552, -71.5833, -96.7541, -106.3833, -110.7333, -112.0167, -108.5333, -93.5781, -118.3667, -84.8948, -95.09, -98.0614, -86.0967, -71.3, -119.3167, -80.55, -100.75, -88.9167, -88.05, -71.4167, -84.23, -75.9833, -80.8536, -101.4, -84.6374, -101.76, -72.0608, -82.4625, -160.8, -100.55, -68.8167, -92.0258, -65.8833, -156.6747, -71.6833, -80.8, -158.0667, -85.1836, -79.3347, -116.5231, -100.9503, -102.1833, -120.12, -83.4764, -78.98, -82.5238, -83.7792, -85.7956, -113.35, -97.6833, -75.6, -98.52, -84.3953, -63.63, -95.32, -124.83, -89.0, -63.4667, -116.1622, -117.1167, -81.4237, -114.4833, -70.8, -79.9, -133.5, -89.2561, -67.38, -105.17, -73.5833, -61.68, -72.52, -76.5501, -98.737, -72.1667, -58.35, -124.4, -77.15, -61.6833, -72.83, -68.15, -118.44, -97.0369, -116.0333, -112.8667, -104.6, -129.9, -125.99, -101.6833, -120.1333, -82.4, -116.1642, -96.2683, -101.5078, -67.1333, -81.1088, -99.3575, -66.6505, -115.55, -121.7667, -59.1667, -93.4389, -131.6, -79.88, -106.9667, -99.2489, -83.6667, -100.0569, -63.52, -81.7667, -82.1794, -104.8483, -140.85, -122.2833, -83.5667, -77.37, -91.15, -79.95, -73.15, -154.3584, -149.65, -96.109, -73.4833, -157.85, -118.0667, -147.62, -147.8667, -113.5103, -112.5006, -85.2333, -64.53, -81.6, -101.8833, -92.88, -80.9486, -98.9327, -88.71, -98.9847, -96.3667, -123.5, -87.68, -81.85, -122.3, -100.5689, -90.68, -88.0667, -119.05, -94.52, -78.6333, -103.6, -152.1, -135.0978, -166.3393, -121.6203, -160.4, -122.6719, -150.1, -95.03, -155.9667, -148.83, -97.8667, -156.0456, -89.8667, -90.2667, -76.5333, -79.4, -77.5333, -81.3833, -85.5833, -99.95, -78.2667, -116.2952, -106.6167, -57.2167, -76.2961, -90.1875, -90.1333, -68.2, -89.2121, -96.75, -71.0, -98.1059, -108.7333, -79.93, -87.781, -76.6, -75.4333, -97.0333, -99.6833, -90.1078, -71.5, -98.4333, -78.38, -117.3333, -106.6167, -78.43, -81.25, -70.708, -122.3833, -102.3167, -83.6, -88.7506, -98.5833, -75.9, -80.8, -128.6442, -94.0667, -88.8486, -120.7333, -98.0799, -89.53, -94.9167, -103.2648, -90.3833, -122.8167, -93.0667, -102.39, -91.5111, -68.3667, -86.75, -83.2, -72.5667, -74.8411, -98.95, -75.3961, -77.9167, -61.8667, -114.8833, -124.4333, -110.2, -94.7, -124.16, -90.4093, -81.7167, -74.6694, -75.85, -97.5667, -84.96, -95.0, -93.22, -96.1833, -79.78, -77.4553, -122.6053, -75.4, -85.1667, -107.2667, -98.6685, -94.73, -88.1167, -100.4086, -67.15, -101.6167, -86.25, -87.6167, -122.4833, -97.7756, -81.75, -162.1104, -102.241, -101.3667, -70.6722, -72.9833, -105.25, -105.048, -63.5167, -75.7167, -103.6833, -91.489, -112.6, -97.3378, -93.8431, -89.3333, -89.6833, -97.4333, -83.44, -100.2856, -80.2329, -94.5, -83.75, -85.5934, -133.35, -84.5208, -58.5661, -64.83, -122.4996, -77.86, -79.03, -70.93, -97.9659, -66.8, -119.65, -100.6, -73.4167, -141.1606, -149.8, -66.4333, -151.25, -164.5, -117.692, -162.0667, -147.0667, -115.1333, -105.1623, -81.6805, -81.3903, -113.5931, -91.5667, -93.032, -95.6567, -70.0667, -84.1889, -159.0499, -94.4014, -81.94, -117.41, -83.0092, -84.5986, -93.3833, -80.7091, -104.6562, -88.8553, -96.1544, -93.5529, -81.33, -83.8333, -73.1667, -93.3, -119.0943, -86.3167, -96.0, -83.4455, -88.2833, -82.8833, -80.2406, -96.7667, -72.8689, -112.1944, -98.6619, -77.7106, -121.25, -94.88, -88.4806, -93.99, -79.851, -95.55, -80.2833, -90.202, -96.6074, 177.57, -76.6667, -86.4333, -98.9565, -92.4516, -86.4, -114.3, -87.4215, -80.2211, -96.3833, -99.75, -121.9333, -78.07, -92.07, -90.6333, -92.91, -86.5, -104.75, -98.891, -117.8086, -75.8655, -85.0525, -97.3496, -81.6833, -98.1211, -75.7, -80.3833, -82.45, -81.1167, -77.95, -90.65, -96.8, -71.12, -116.6167, -96.43, -95.8633, -87.1668, -93.25, -106.72, -71.1739, -81.97, -113.7661, -159.35, -91.4156, -73.75, -137.2333, -99.84, -78.8333, -78.74, -105.62, -81.74, -97.6, -117.3494, -93.3269, -95.95, -86.059, -78.15, -121.4, -90.4722, -120.5139, -84.63, -82.5, -94.7167, -100.5833, -95.395, -92.1407, -81.3167, -83.65, -83.7374, -86.2833, -107.9, -82.2667, -93.3833, -97.0972, -103.2008, -110.7333, -80.2333, -102.6525, -115.6734, -119.3, -67.25, -63.5667, -99.3381, -99.0, -121.2367, -64.6833, -80.3, -98.2167, -112.0167, -62.6833, -81.4236, -76.4944, -122.2208, -106.0095, -75.25, -82.5289, -74.53, -133.05, -119.2833, -118.32, -116.5, -116.47, -66.25, -115.78, -109.5, -92.6912, -123.2667, -99.2667, -71.27, -123.47, -138.9167, -71.22, -80.6167, -105.93, -112.67, -90.4667, -114.2192, -123.2333, -72.7875, -54.8, -59.63, -82.4167, -113.6333, -57.58, -107.9558, -89.65, -74.6, -117.0903, -112.8167, -123.43, -97.4167, -96.943, -80.55, -124.4667, -82.4493, -115.5753, -113.95, -87.9833, -98.32, -88.4667, -71.03, -115.0667, -89.7, -80.6344, -76.0264, -97.7953, -84.9, -113.889, -72.885, -111.45, -96.15, -91.98, -84.05, -91.88, -90.9167, -84.8, -75.6667, -84.5667, -106.9475, -70.9167, -91.65, -98.9, -84.7697, -122.4208, -114.8611, -80.4, -96.0, -98.0558, -112.0656, -89.4076, -95.7826, -95.6667, -149.45, -72.5369, -82.1547, -122.5833, -88.1333, -98.3167, -97.8333, -85.5167, -70.5333 ;
       station_name = "CYFC", "K9MN", "KDDC", "KVQQ", "KDDH" ; //, "KOTM", "PAZK", "KOTH", "KOTG", "KBXK", "CYVV", "CYVR", "CTZE", "CYVQ", "K3LF", "MUCU", "KVNY", "CTZR", "CYVC", "MUCM", "MUCL", "CYVO", "KNHK", "PADE", "CYQF", "CYDQ", "PADK", "PADM", "PADL", "KTVL", "PADQ", "PADU", "CYDN", "CXTH", "KOXV", "CYDB", "KPAH", "CYDF", "PPIZ", "KFPK", "KADM", "KO54", "KPAN", "KADC", "KW99", "KADF", "KADG", "KSDB", "KSDA", "KLLQ", "KFPR", "KADS", "KADU", "KSDL", "KADW", "KMRF", "KMRB", "KMRN", "KMRJ", "KMRH", "KMRT", "KMRY", "KTVI", "PHMK", "KSRC", "KSRQ", "KSRR", "KRCE", "KJBR", "KVCV", "KVCT", "KOZW", "KBJI", "KOZR", "KBJJ", "KRCX", "KBJC", "KVCB", "KOZA", "KWST", "K2WX", "CWEQ", "CWEP", "CWEW", "CWEI", "CWEH", "CWEK", "CZKA", "K11R", "CWEO", "CWEA", "CWEC", "CWEB", "CWFJ", "CXKM", "KTOP", "KTOR", "CXKE", "CXKA", "KTOA", "KTOB", "KTOL", "KTOI", "KTAZ", "KMLT", "KMLU", "KMLP", "K06D", "KTAN", "KMLI", "KMLJ", "KMLE", "KTAD", "TJSJ", "KMLB", "KMLC", "KGOP", "KGOV", "KDYR", "K2C8", "KIOW", "KGOK", "KGON", "KBDL", "KRQO", "KFHB", "KRQE", "KRQB", "KEKQ", "KGSB", "KGSO", "KGSH", "KSMX", "KNYL", "KGSP", "KNYC", "KAKO", "KEKO", "KNYG", "KROG", "KROC", "KPOV", "KROA", "KEYW", "KROW", "KPOB", "KPOE", "KPOF", "K08D", "KEYF", "KEYE", "KWAL", "KHGR", "CYFS", "CWKP", "CWKX", "CWKG", "CXYH", "CWKB", "CWKO", "CYDL", "CWKM", "KRAP", "KPSF", "PAKI", "PAKK", "KPSM", "KPSN", "KPSO", "KLPC", "KNKX", "CYET", "CYEK", "KPSP", "CYEN", "CTKG", "PAKT", "PAKU", "PAKV", "PAKW", "KPSX", "CYED", "KFSW", "KFST", "KJSV", "KIPT", "KJST", "KAEL", "KSET", "KFHU", "KAEG", "KSEP", "KSHV", "KLKR", "KAEX", "KLKU", "KLKV", "KFSO", "KSEG", "KFSM", "KSEA", "KJSO", "KFSI", "KCKC", "KADH", "KHUL", "KHUM", "CWYI", "KASX", "CWYJ", "KHUF", "KAST", "KCKI", "KFAT", "KCKN", "KCKM", "KHUA", "KCKP", "CWYY", "KCKV", "KASJ", "KASE", "KASD", "KHUT", "KUGN", "CWYQ", "KFAF", "KDUJ", "KSHN", "KDUH", "KDUC", "KDUA", "KDUG", "KDUX", "CWZW", "KXVG", "CWZQ", "KSSI", "KSDY", "KSSC", "K5H4", "CWZS", "KSSF", "KJEF", "PFNO", "KJER", "KJES", "CPQW", "KBMI", "KVBS", "KBML", "KVBT", "KONO", "KBMG", "KVBG", "KSDF", "KVPZ", "KVPS", "KDCM", "KDCU", "KOUN", "KVPC", "PAYA", "K3MW", "CYMM", "KONZ", "PHNY", "CYWA", "PHNG", "CYWG", "CYWK", "KSDM", "CYWL", "KKLS", "KCEF", "CWJH", "KMMV", "KMMU", "KMMT", "KMZZ", "KMML", "KMMK", "KMMH", "KLWD", "KGLY", "KGLW", "KGLR", "KGLS", "KGLH", "KCEY", "KGLD", "KGLE", "CTWL", "KCEZ", "KMSL", "KMSO", "KMSN", "KMSP", "KMSS", "KMSV", "KMSY", "K1U7", "PAFE", "KPNS", "KRND", "KPNT", "KRNH", "KRNM", "KRNO", "KPNC", "KRNP", "KPNA", "KGBG", "KRNT", "KPNE", "KGBN", "KPNM", "KGBK", "KEZF", "CWHP", "CWHQ", "CWHV", "CWHT", "CAMS", "KCZZ", "KEZS", "KCKB", "KHFD", "KHFJ", "CWHN", "CWHL", "CWHM", "K12N", "KTNU", "KIRS", "K8A0", "KTNX", "KIRK", "KTNB", "KHIF", "KATY", "KMER", "KHTL", "KATP", "KCHD", "KATS", "KATT", "KCHA", "KATL", "KIFP", "KHTS", "KCHS", "KDTW", "KTPA", "KDTS", "KNUQ", "KDTL", "KDTO", "KDTN", "KRPJ", "KRPH", "KRPD", "KNXX", "KEDU", "KGPI", "KGPM", "KECU", "KCAO", "KGPT", "GA45", "KGPZ", "KEDE", "KRWL", "KNXF", "KEDC", "KT82", "KAWM", "CVTS", "KDBN", "KDBQ", "KBZN", "KVSF", "CYXX", "CYXY", "CYXT", "CYXU", "CYXP", "CYXR", "CYXS", "CYXL", "CYXH", "PHOG", "CYXD", "CYXE", "CYXC", "KPRG", "PAJN", "KPRC", "KPRB", "K3J7", "KPRO", "KPRN", "PAJC", "KPRS", "PAJZ", "KNJK", "KNJM", "KPRX", "PFYU", "KAFW", "KHZE", "CWVF", "KAFP", "KSBP", "KSBS", "KAFF", "KCFV", "KSBM", "KFRG", "KSBO", "KAFN", "KSBA", "CWZV", "KFRM", "KAFK", "KHZY", "KHZX", "PATQ", "KP69", "KP68", "KP60", "CWVQ", "CWVT", "CWVU", "KSPW", "KSPR", "KSPS", "KJDD", "KSPF", "KSPG", "KSPD", "KBJN", "KSPB", "KSPA", "KSPI", "KOXR", "KBLI", "KBLH", "KL63", "KBLM", "KBLF", "KOXB", "KOXC", "CWWK", "KOXI", "KBLV", "KBLU", "K1V4", "PATC", "CZMJ", "CZMD", "CXIB", "KTMB", "KISM", "KTMA", "CMMY", "KTME", "KTMK", "KMNZ", "KONL", "KONM", "K04W", "K04V", "KONA", "KONX", "KMNH", "KMNI", "KMNN", "KMNM", "KONP", "K0J4", "KONT", "KMNE", "K2J9", "KIAH", "KIAG", "KIAD", "KGMU", "KIAB", "KGMJ", "KGCC", "KXNA", "KRDR", "KE80", "MDPC", "KRSP", "KRSV", "KRSW", "KRST", "CWEZ", "KRSN", "KRSL", "KGCM", "KGCK", "KEET", "KPCZ", "KEEO", "KEEN", "KPCM", "KEED", "KRAL", "KTTD", "KPMV", "KISO", "KISN", "KPMP", "KRAC", "KISW", "KGCD", "KISQ", "KISP", "KGCN", "KPMD", "CNVQ", "KRAS", "CWIY", "CWIX", "CWIZ", "CWIT", "CWIW", "CWIS", "KHEQ", "CWIL", "CWII", "CWIK", "KHEI", "KHEF", "CWEL", "PAIK", "PAII", "PAIN", "PAIL", "PAIM", "KPQI", "KPQN", "PAIG", "KPQL", "KNEL", "KPHP", "CYKA", "PAIW", "KCGF", "KAGS", "KAGR", "KCGC", "CYBU", "KLIC", "KCGI", "CYGQ", "KHYS", "KAGC", "KSCH", "KCGS", "KHYW", "CYGW", "CYGV", "CYGX", "KLIT", "KCGZ", "KCIN", "KAUS", "KCIC", "KAUW", "KCID", "CAPR", "KAUH", "KAUO", "KHKA", "KAUM", "KCIR", "KCIU", "KDSV", "KFCM", "KFCI", "KFCS", "TNCM", "TNCC", "TNCB", "TNCA", "KDSM", "TNCE", "KLGD", "KLGA", "KLGB", "KLGC", "KJGG", "KSQI", "KSJT", "K7L2", "KSQL", "KNGU", "KBOW", "KSAZ", "KBOS", "KLNC", "KCCR", "KDOV", "KVLL", "CXSR", "KVLD", "KBOK", "KBOI", "KDAN", "KDAL", "KNEW", "KP53", "KW22", "KDAG", "KDAB", "KW29", "KP58", "KP59", "CXKT", "KZZV", "KDAY", "KDAW", "CTGT", "KVRB", "CYYZ", "CYYY", "CYYU", "CYYR", "CYYQ", "CYYN", "CYYL", "CYYJ", "CYYG", "CYYF", "CYYE", "CYYD", "CYYC", "CYYB", "KOOA", "KUVA", "KDZB", "KMOD", "KMOB", "KMOT", "KMOP", "CVSL", "KMOX", "KDFI", "K7BM", "KCGE", "KHYA", "KMLS", "KABY", "CWTS", "KHYI", "KITH", "KPLU", "CYGL", "KITR", "KPLN", "KAJG", "KMLF", "KHYR", "CWNZ", "KETH", "CYGP", "CWNP", "CWNQ", "KETB", "KETC", "CWNH", "KWDG", "CWNK", "CWNM", "KHDO", "KHDN", "KHDC", "CWNC", "KHDE", "CWNE", "K14Y", "KWVL", "KHYX", "CXHR", "KI16", "KSCF", "TAPA", "CXHA", "KTLH", "CXHM", "CXHI", "MKJS", "MKJP", "CAQY", "KCVS", "KLZZ", "KCVX", "KCVG", "KCVB", "KHJO", "KCVN", "KCVO", "KCVH", "KHJH", "KAVC", "KFBG", "KDRT", "KAVL", "KHKS", "KFBL", "KDRA", "KAVP", "KDRI", "KDRO", "KF05", "KIDP", "KDVO", "CAOH", "KHKY", "CAOS", "KTZR", "KDVN", "KHVS", "KGVL", "KRRL", "KEFT", "KPBX", "KGVX", "KRRT", "KGVT", "KEFD", "KAUN", "KHVR", "KT65", "KFVE", "CYZX", "CYZY", "CYZR", "KUAO", "CYZP", "CYZV", "CYZT", "CWPR", "CYZH", "KHNR", "KDLS", "CYZE", "KPPO", "KN60", "KPPF", "KPPA", "PAKN", "PAHC", "PAHL", "PAHO", "PAHN", "KPPQ", "KCDC", "KCDA", "KLHM", "KCDD", "CYHK", "CYHD", "CYHE", "KCDH", "KLHB", "KCDN", "KAHQ", "K9A1", "KCDR", "KCDS", "KAHN", "KLHZ", "KCDW", "KY19", "KCNU", "KLHQ", "KULM", "KLHW", "KBPT", "KENL", "CTTR", "KCNM", "KEBS", "CYNM", "KENV", "KHND", "K4BM", "KCNI", "KJFX", "KJFZ", "KLFK", "KLFI", "KLFT", "K1F0", "KJFK", "PASK", "KACV", "KBNW", "KDNN", "CERM", "KDNK", "KNBT", "KBNA", "KDNV", "KDNS", "KLRD", "KBNL", "KBNO", "KWWR", "CXVN", "K3T5", "KWWD", "CZOC", "CXOX", "CXOY", "KTKV", "KTKI", "KTKC", "KOLV", "KOLU", "KOLS", "KOLZ", "KOLY", "KOLF", "KOLE", "KOLM", "KICT", "KMHE", "KLGU", "KMHK", "KRDD", "KMHR", "KMHS", "KMHT", "KMHV", "KICL", "KEKN", "KTYR", "KTYS", "KTYQ", "KBHK", "KPOU", "KGWO", "KRUE", "KRUG", "KGWB", "KRUQ", "KSWW", "KRUT", "CWYL", "KPAE", "KD50", "CYIV", "KGWW", "KPAO", "KD55", "CNPK", "KRCM", "KRCA", "KTVR", "KRCZ", "KGAO", "KGAI", "KRCR", "KGAD", "KGAG", "KGAF", "CWOY", "KEUL", "KEUG", "KEUF", "KCYS", "CWOV", "CWOK", "CWOI", "CXBD", "CWON", "KYIP", "CWOC", "CWOE", "CWOD", "PAOR", "KPWK", "PAOT", "PAOU", "KPWA", "KNGP", "KPWC", "KPWG", "CWBT", "KTVF", "PAOH", "KPWT", "PAOM", "PAOO", "KLWT", "KLWV", "KAIZ", "KLWS", "KTVC", "KAIT", "KCEC", "KAIO", "KAIK", "KLWA", "KLWB", "KLWC", "KAIG", "KLWM", "KCEW", "KAID", "KWMC", "KAIA", "KEGE", "KCWV", "KNUI", "KLYV", "KUCP", "CARP", "KEGI", "KHIB", "KCWF", "KEGV", "KCWC", "KCWA", "KHIE", "KNUW", "KHIO", "KCWI", "KFMN", "KFMH", "KAWG", "CXSC", "KFME", "CXSH", "KAWO", "KLYH", "KFMY", "KDQH", "KLEB", "KLEE", "K3I2", "KLEW", "KRBL", "KLEX", "KHXD", "KDMA", "KBAX", "KBAZ", "KDMH", "KDMN", "KDMO", "KEFK", "KDMW", "KBAD", "KBAF", "KCMY", "KBAB", "MDPP", "KJWG", "KSAC", "KSAD", "KSAF", "KSAN", "KSAR", "KSAT", "KSAW", "KSAV", "KDAA", "KO22", "KJWY", "KCEU", "PHBK", "CVQZ", "K4A9", "CTKR", "KOMA", "KOMH", "KOMK", "KMIC", "KMIB", "KMIA", "KJXI", "KMIE", "KPSC", "KL35", "KIDA", "KMIW", "KMIV", "CYER", "KIDI", "PAKF", "PASD", "PASA", "KVNC", "PASC", "PASL", "PASM", "PASN", "PASO", "PASH", "PASI", "CYEV", "PASV", "CWPU", "KVNP", "KPSK", "PASX", "PASY", "PAKP", "CZPC", "KRBW", "KLOT", "KRBD", "KRBG", "KGFK", "KGFL", "KGFA", "KRBO", "KMBS", "K4O4", "KEVM", "CYEG", "CACP", "CZPK", "KWJF", "KEVV", "KEVW", "CPIF", "CPIL", "K36U", "PABT", "KI39", "CXNP", "KSHD", "KSEZ", "KTCC", "KHSI", "CXNM", "CWRY", "CWRZ", "KCTZ", "CWRU", "CWRV", "KCTY", "KLXT", "CWRR", "KHHR", "KCTB", "CWRM", "CWRN", "CWRO", "CWRH", "KLXL", "CWRJ", "KLXN", "KCTJ", "KNTU", "KHHF", "KFLO", "KAXN", "KFLL", "KAXH", "KFLG", "KFLD", "KAPG", "KAXA", "KPBH", "KFSE", "KAXX", "KDPL", "KFLY", "KDPA", "KFLP", "CWLF", "CWLE", "CWLB", "CWLC", "CWLM", "CWLJ", "CWLI", "CWLV", "CWLS", "CWLP", "KTXK", "CWLY", "KIXD", "KGTU", "KGTR", "KIXA", "KRTN", "KGTF", "KGTB", "KSNL", "KFAY", "KSBY", "KSNA", "KSNC", "KSNY", "KSNT", "KSNS", "KNBG", "CWYE", "KPBF", "KFAR", "KPVJ", "PANW", "PANV", "PANT", "KPVC", "KPVB", "KPVG", "KPVD", "PANC", "PANI", "KPVW", "PANN", "KPVU", "KNFE", "KSHL", "KNFG", "KCBK", "KUNV", "KWYS", "KUNU", "KNFL", "KIBM", "KCBE", "KCBF", "KCBG", "KNFW", "KASN", "KAJO", "CWPG", "KLVN", "KLVM", "KUNI", "KLVK", "KUNO", "KNSI", "KFAM", "PARC", "KVIH", "CTRA", "KVIS", "PARS", "KMXF", "KASG", "PARY", "KMXO", "CWWE", "CWRT", "CWPE", "KCNO", "CMFM", "KLDM", "KNTD", "KUXL", "KJHW", "KLXV", "K1H2", "KDLL", "KDLN", "KXMR", "KDLH", "K42J", "KDLF", "MDSD", "KDLZ", "K7A7", "MDST", "CWRK", "CWRD", "CXMW", "KROS", "CXMP", "CXMM", "CXMI", "CXMD", "CXRG", "KOBE", "KIER", "KIEN", "KMJQ", "CTPQ", "CWME", "CWMI", "CWMJ", "CWMM", "KBBG", "CWMQ", "KTWM", "PAPN", "CXCA", "CABR", "CWMX", "K8D3", "CXRH", "CABT", "CXCK", "KGUP", "KGUS", "KRWI", "KRWF", "KD39", "KPGV", "KGUC", "KRWV", "KPGA", "KPGD", "PAPG", "KIWI", "KIWA", "KMDH", "KTIK", "KMDJ", "KMDT", "KTIW", "KNKT", "KMDW", "KRXE", "KMDQ", "KTIP", "KMDS", "PAPB", "KGGG", "KMDZ", "KREO", "KYKM", "KYKN", "KEWR", "CZSP", "CZSJ", "KUBE", "KEWB", "KEWN", "KEWK", "KPUW", "CVAS", "CMTH", "PAMY", "PAMR", "KRYT", "PAMO", "KRYV", "PAMM", "KPUB", "KPUC", "PAMH", "PAMD", "KPUJ", "PAMC", "KCNC", "KCCO", "KUOX", "KLUX", "KNAK", "CYKY", "CYKZ", "KCCY", "KEDW", "KLUF", "KLUD", "KLUK", "KCCU", "KLUM", "CWSY", "KHOP", "KCUT", "CWSU", "CWST", "KHOT", "KHOU", "CWSP", "KCUL", "CWSL", "CWSK", "KCUH", "KEAU", "KEAT", "CWSG", "CWSF", "KHOB", "CWSD", "KHOE", "CWSA", "KCUB", "KFOK", "KFOA", "KFKN", "KFOD", "KFOE", "KFOZ", "KAYS", "KLCH", "KLCI", "KLCK", "KLCG", "KJKJ", "KJKL", "K9D7", "KJKA", "KDKK", "KDKB", "KBCT", "KBCK", "KBCB", "KDKR", "KXLL", "KBCE", "KJYL", "KJYM", "KJYO", "KP92", "KFYJ", "KJYG", "KAKH", "KSOA", "KAKQ", "KFYV", "KAKR", "KSOW", "KJYR", "KSOP", "KMGR", "PACV", "KBQK", "PACZ", "PACD", "PACM", "KBQP", "K1P1", "KDCA", "KOCW", "KDXX", "KOCH", "KOCF", "KMKJ", "KMKL", "KMKO", "KMKN", "KMKC", "CWVO", "KMKE", "KMKG", "KMKS", "KMKT", "KIFA", "KMYR", "KMYP", "KMYV", "KMYT", "KMYF", "PAQT", "KWDR", "KMYL", "KCXY", "KHEZ", "KC09", "KHBR", "KAUG", "KMEB", "KRDU", "KMEM", "KMEI", "KMEH", "KRDG", "KCXP", "KTHV", "KRDK", "KMEZ", "KRDM", "KGDB", "KCXO", "K4M9", "KGDJ", "KGDV", "KGDP", "KEPH", "K4MR", "KJVL", "CPOX", "KLMT", "MUVR", "KLNP", "CXLT", "CXLL", "KCLS", "CXLB", "CWPZ", "KHNZ", "CWPX", "KCRP", "KCRQ", "KCRS", "KCRW", "CWPK", "CWPN", "CWPO", "CWPL", "KHNB", "CWPF", "KCRE", "CWPD", "KCRG", "KFNT", "KAZO", "CXPA", "KFNB", "KFNL", "K96D", "CXPS", "CWBM", "KC75", "CWBO", "CACQ", "CXBR", "CXBQ", "CWBK", "CWBD", "CWBE", "CWBA", "CWXR", "MMSP", "KTVK", "CWBY", "CWBZ", "CXBO", "CWBU", "CWBV", "CXBK", "PHNL", "CXBI", "CWBS", "KIZA", "KIZG", "KWVI", "KGZL", "KGZH", "KRVS", "KJXN", "KALB", "KSLI", "KSLN", "KSLO", "KFXE", "TJPS", "KSLB", "KALI", "KALK", "KALM", "KALN", "KALO", "KALS", "KALW", "KALX", "KFXY", "KACB", "PABV", "KVYS", "KBPK", "PABR", "KBPI", "CMGB", "KBPG", "KBPC", "KDEH", "CTBT", "PABE", "PABA", "PAHY", "KACY", "PABL", "PABI", "KPTS", "KPTT", "KPTW", "KPTV", "PALP", "PALU", "PALH", "KPTB", "KACT", "KPTK", "PALG", "KPTN", "KELD", "KY51", "KY50", "CYLW", "KELM", "KELN", "KELO", "KLTS", "KACP", "PHSF", "KELP", "CYLH", "CYLL", "KELY", "KELZ", "KORL", "KBBD", "PAPO", "KBBF", "KORH", "PAPH", "KBBB", "KORD", "KORE", "KORF", "KORG", "KORB", "KORC", "KBBW", "KMZJ", "KBBP", "KMZH", "KVKY", "KMZG", "KRGK", "KORS", "CYPD", "CYPE", "CYPA", "CYPH", "CYPQ", "CYPR", "KCHK", "CYPY", "KLBL", "KLBB", "KLBF", "KLBE", "KLBX", "KUZA", "KLBR", "KLBT", "K40J", "KHSB", "KSZL", "KSZT", "KMDD", "KLZU", "KUES", "CZCR", "CZCP", "KLVS", "KCBM", "KIGX", "KMTV", "KMTW", "KMTP", "KVEL", "KIGM", "KVER", "KMTC", "KMTN", "KMTO", "KMTH", "KMTJ", "CWCO", "CZUB", "CWCL", "CWCJ", "CWCH", "CWCF", "KTUP", "CZUM", "CWCA", "KNZY", "CXAF", "KTUL", "CWCT", "KRIV", "KRIW", "KDRM", "KSLK", "KRIC", "KRIL", "KHQZ", "KASW", "KMFD", "KMFE", "KMFI", "KIIY", "KMFR", "KSLH", "KMFV", "KIIB", "KGED", "KGEG", "KEQY", "KLVJ", "KROX", "K6R3", "KFSD", "KGEU", "CYJT", "K6R6", "KGEY", "KGEZ", "KAVK", "KCOQ", "KCAR", "CYMT", "KHST", "KHSV", "CYMX", "KHSP", "KLSV", "KNCA", "KEMV", "CYMA", "KCAE", "KUIN", "KCAG", "KUIL", "KHSE", "KCAK", "CYMO", "KLSE", "KLSF", "PHTO", "KPEF", "KPEA", "KNQX", "KPEO", "KCSQ", "KCSV", "KECG", "KNQA", "KCSM", "KPEQ", "KNQI", "KCSG", "KPEX", "CWQD", "KFIT", "CXWM", "CXWN", "KHMN", "CWQL", "CWQH", "CXWF", "KIGQ", "CWQW", "CWQV", "CWQQ", "KAVX", "CWQS", "KFIG", "KLAW", "KLAR", "KLAS", "KNMM", "KLAX", "KLAF", "KLAA", "KLAN", "MUHG", "KLAL", "KLAM", "MUHA", "KSLC", "KFUL", "KY63", "KXBP", "KJMR", "KJMS", "KDIJ", "KDIK", "KAMA", "KAMG", "KSMP", "KSMS", "KBMQ", "KVES", "KAMN", "KSME", "KSMF", "KAMW", "KSMO", "KSMN", "PAAQ", "KOEO", "PAAK", "KLLJ", "KASH", "K21D", "KSLG", "KVDF", "KMUT", "KPWM", "KVDI", "KOAJ", "KTUS", "KMUO", "KMUI", "KVJI", "PAWI", "KBED", "PAWN", "KOSH", "KBEH", "KOSC", "CWWA", "KOSA", "PAWG", "KCQB", "KSLE", "KOSU", "PAWS", "K9L2", "CYQG", "KGBD", "CYQD", "CYQB", "CYQA", "CYQM", "CYQL", "CYQK", "PHHI", "CYQI", "CYQH", "CYQW", "CYQV", "CYQU", "CYQT", "TIST", "CYQR", "CYQQ", "TISX", "KHWD", "CYQZ", "CYQY", "KMGM", "KMGN", "KMGJ", "KMGE", "K0VG", "KIJX", "KFKS", "KRFI", "TJNR", "KMGY", "KIJD", "KMGW", "KRFD", "KTFP", "KEBG", "KPBG", "KERY", "KERV", "KYNG", "KERI", "KGJT", "KIPJ", "CWWZ", "KI75", "KD07", "CZBF", "KPBI", "CAHK", "KPDC", "KPDK", "KNPA", "KPDT", "KPDX", "KFHR", "KHLC", "CWVC", "KCPC", "KHLG", "CWVI", "K0A9", "CXVG", "KCPK", "CWVN", "KHLN", "CWVP", "KCPW", "KCPT", "KHLR", "KCPR", "KCPS", "KHLX", "CAWR", "KHFF", "CZTB", "KRHV", "KGXY", "KTTA", "KSLR", "KRHP", "KTTN", "KSIY", "KTTS", "KRHI", "KSJS", "KANJ", "KANK", "KSJX", "KAND", "KANE", "KANB", "KFZG", "KFZY", "KSJC", "KFFX", "KANW", "KJZI", "KSJN", "KXSA", "CVLY", "KBRD", "CYUX", "KBRL", "KBRO", "KRZL", "KRZN", "KAAF", "KPZQ", "KHPN", "CVBB", "KCNY", "KEND", "KHRX", "KY70", "KNBC", "KHRT", "KLRU", "KHRO", "KLRJ", "KHRL", "KLRO", "KENW", "KHRI", "KCNK", "CYNE", "KLRF", "KCNB", "CYNA", "KOPN", "KBDE", "PAVL", "PAVC", "PAVA", "KBDH", "KOPF", "KBDN", "PAVD", "KBDR", "CBBC", "KBDU", "KVUO", "KGGI", "KVUJ", "CYRJ", "PHIK", "CYRV", "CYRT", "MUGM", "K2G4", "KNLC", "KUTS", "KUTA", "KFTG", "KDHT", "KNDZ", "KFTN", "KFTK", "KJLN", "KDNL", "KFTW", "KSXT", "KFTY", "KDHN", "PALJ", "K33V", "PAHP", "KM19", "CVOD", "CZEV", "CZEL", "KSKX", "KSVC", "K20V", "KSVN", "KGEV", "KSVH", "K1A5", "MYNN", "KOFF", "KMVY", "KOFP", "KVGT", "KMVE", "KMVN", "KMVL", "KSKF", "CZWN", "CWAV", "CWAQ", "CWAS", "KCHO", "KAQR", "CXGH", "CWAF", "CXGM", "CAFC", "CWAJ", "KRKR", "KRKS", "KRKP", "KGNA", "KTSP", "KRKD", "CYHM", "KTEB", "KIKW", "KIKV", "CVOP", "KIKR", "KTEX", "KIKK", "KATW", "KTEW", "KGKJ", "KEST", "KCDJ", "KGKY", "KESN", "KESC", "KESF", "KC29", "KPYX", "KGGE", "KPYM", "CYOY", "KEOK", "KLHX", "KEOE", "KCOU", "KCOT", "KCOS", "CYOW", "KHQU", "KCON", "KCOM", "KHQI", "CYOO", "KHQM", "KCOF", "KCOE", "KCOD", "CYOD", "KDYS", "PAGN", "KGYB", "KPKD", "KGYL", "KGYI", "KGYH", "KPKB", "KGYR", "KPKV", "KNSE", "KGYY", "CWWC", "CWWB", "KCQC", "CAHW", "CWWF", "CAHR", "K9V9", "KHCD", "KCAV", "KCQM", "CWWN", "CWWL", "CAHD", "KFKL", "CWWP", "KCQT", "KCQW", "KGNR", "KCQX", "KFKA", "KNOG", "KLOZ", "K5C1", "KLOU", "KUUU", "KLOR", "KLOL", "KLOM", "CYAM", "CYAH", "KFWC", "KFWA", "KSYM", "KAAA", "KSYN", "KAAO", "KDGW", "KFWN", "KFWS", "KPIE", "KAAT", "KJOT", "KSYR", "KCAD", "KFET", "KAOH", "KFEW", "KFEP", "KAOO", "KUKF", "KUKI", "KEMP", "KLQK", "KSKA", "KUKT", "PAGY", "KBUR", "CVOQ", "KDYB", "KBUU", "CVOU", "KBUY", "KDYL", "PAGS", "PAGH", "CVOC", "KDYT", "PAGK", "PAGL", "PAGM", "KBUF", "PAGA", "CVOI", "CVOM", "KSWF", "K1M4", "KSWO", "KJAN", "K3A1", "KJAS", "KJAX", "KS25", "KBID", "KBIE", "KBIF", "KJAC", "KOGD", "KBIL", "KMWT", "KBIH", "KBIJ", "KMWM", "KMWL", "KBIV", "KMWN", "KMWH", "KMWK", "KBIS", "KBIX", "KMWC", "KOQU", "KOQT", "KBGM", "KOGB", "KBGD", "KBGE", "KOGA", "CMLU", "KVTA", "PAUN", "KVTN", "KBGR", "KVTI", "CYSJ", "PHJH", "CYSC", "CYSB", "PHJR", "KMAI", "KMAO", "KMAN", "KSNK", "KMAF", "KMAE", "KTDZ", "KTDF", "K4I3", "KILN", "KECP", "CXCP", "KILE", "KILG", "KPEZ", "KMWO", "CABB", "KGHW", "CWQC", "KMWA", "CZDB", "KNXP", "KNRS", "KNRB", "KTWF", "CWTN", "KHBI", "CXTV", "KHBG", "CWTG", "KVTP", "CWTA", "CXTD", "CWTY", "K2W6", "KHBV", "CWTT", "CWTU", "CXTL", "CWQP", "CWFP", "CWFQ", "CWFW", "CXFR", "KWLD", "CXFV", "CWFE", "CWFF", "CWFG", "CXFA", "CWFO", "KTRK", "KTRI", "KTRM", "KTRL", "KGUY", "TJBQ", "KFDW", "CWZE", "CWZF", "CWZG", "CWZA", "CWZB", "CTAG", "CWZL", "KUDG", "KSHR", "KAPY", "KFDY", "CWZT", "CWZU", "KAPF", "KLPR", "KAPA", "CWZR", "KAPC", "KAPN", "KFDK", "KBTR", "KBTP", "KBTV", "PAFS", "PAFR", "KBTA", "KDXR", "PAFM", "KMWS", "PAFB", "PAFA", "KDXZ", "KBTM", "KBTL", "TUPJ", "KEHO", "KEHA", "KEHC", "KCLT", "KCLK", "KCLI", "KFDR", "KCLL", "KCLM", "KEHR", "KCLE", "KBFI", "KTIF", "KOVS", "KBFM", "KBFL", "KVWU", "KBFD", "KBFF", "PATA", "CVXY", "PATE", "KOVE", "PATG", "CVXS", "PATK", "KOVL", "PATL", "PATO", "CYTH", "PHKO", "CYTL", "KVOK", "CYTE", "CYTZ", "CYTR", "CYTS", "KPAM", "CYBR", "CTNK", "K65S", "KGGW", "CYBX", "KLNS", "KLNR", "KIWD", "CYBC", "KLNL", "KLNK", "CYBG", "KS32", "KLND", "CYBN", "KVOA", "KSFQ", "KABE", "KDFW", "KABI", "KSFY", "KSFZ", "KABR", "KJNX", "KSFF", "KABQ", "KFVX", "KSFB", "KSFM", "KSFO", "CZHB", "KWRB", "KM30", "KP28", "K2DP", "KTIX", "CZGH", "KSTC", "KSTF", "CYXJ", "K2D5", "KSTE", "KSTJ", "KSTK", "KSTL", "KSTS", "KSTP", "KODO", "KMPZ", "KBHB", "KBHM", "KVAD", "KMPV", "KVAY", "KODX", "KMPO", "KILM", "CWGR", "CWGW", "CWGT", "CWGY", "CWGX", "CWGB", "K1R7", "CWGD", "KSMQ", "CWGH", "CWGN", "KRMY", "KTQH", "CXEA", "KTQE", "CXET", "KRMN", "KO69", "KRME", "KRMG", "KTCS", "KOJA", "KOJC", "KIMT", "KMBG", "TJMZ", "KIML", "KMBL", "KTCL", "KTCM", "K0F2", "KGIF", "PAMK", "K2V5", "CWXB", "KGHG", "CMRF", "CWXG", "KEIK", "CYHZ", "CXOA", "KE38", "KEIR", "KPIH", "KPIL", "KCFE", "KPIB", "KPIA", "KOFK", "KTTF", "KPIR", "KPIT", "KLJF", "KARB", "KHAI", "CWUM", "KHAO", "CAJT", "CWXS", "KHAF", "KCJR", "CWUY", "CWUX", "KRYW", "CWUP", "CWUS", "CWUT", "CYHU", "PAEG", "PAED", "CYCX", "PAEN", "PAEM", "KNID", "PAEH", "PAEI", "CYCO", "KLMO", "KNIP", "CTMS", "KSGU", "KSGT", "KSGS", "KSGR", "KACK", "KACJ", "PAMB", "KDEQ", "KFQD", "KDEW", "KDET", "KRYY", "KSGF", "KJQF", "KDEN", "KDEC", "KARM", "KACQ", "KSGJ", "KSGH", "KAQW", "KAQV", "KCMA", "KSBN", "KAQP", "KCFS", "KCMI", "KCMH", "KHWO", "KFRI", "KHWV", "KCMR", "KAQO", "KHWY", "KSCK", "KFGN", "KCMX", "KMGG", "KSIF", "KDWH", "KAFJ", "KXPY", "KBWP", "UHMA", "KBWI", "KBWG", "KBWD", "KCCA", "K79J", "KSUN", "KSUE", "KSUA", "KSUX", "KJCT", "KSUU", "KSUT", "KSUW", "KSUS", "KBKB", "KMQY", "KBKF", "KBKD", "KBKE", "KMQS", "KOEB", "KBKN", "KBKL", "KBKS", "KMQI", "CYKF", "KBKV", "KBKW", "KBKT", "KMQB", "KBKX", "KMQE", "KBYS", "KVVV", "KBYY", "KOWB", "KOWA", "KBYG", "KOWD", "KVVG", "KBYI", "PHLI", "KBFW", "CYUL", "CYUA", "KICR", "CYUY", "KHRJ", "CYKJ", "KTBR", "KOKC", "KOKB", "KMCW", "KOKM", "KOKK", "KOKV", "KMCC", "KMCB", "KMCE", "KMCD", "KMCF", "KMCI", "KMCK", "KMCJ", "KTBN", "KMCO", "KMCN", "K1A6", "KIND", "KGNT", "KGNV", "KINL", "KINJ", "KINK", "KINW", "KINT", "KGNC", "KINS", "CWSV", "CWSS", "CWSR", "KAXS", "KEAR", "CZFS", "TXKF", "KEXX", "KHON", "KPHX", "TKPK", "KPHD", "KPHF", "KOAK", "K0E0", "KPHL", "KPHN", "CWJT", "CWJU", "CWJV", "CWJW", "CWJR", "CZZJ", "CXZV", "CXZU", "CWJX", "KH21", "CWSB", "CWJD", "CWJB", "CWJL", "CWJN", "CWJO", "CXZC", "CWJI", "CWDZ", "CWDV", "CWDU", "CWDR", "CWDQ", "CWDO", "CWDM", "CWDJ", "CWDK", "CWDH", "KWRL", "MMMD", "KWRI", "KTPH", "CXDB", "CXDE", "KTPL", "KHCO", "CXDI", "CXDK", "KTPF", "KIPL", "CXDP", "KIPN", "CXDW", "KARR", "CWXC", "CWXA", "KARV", "KARW", "KART", "KBEA", "KFFT", "CWXN", "KHVN", "CWXL", "KFFM", "KFFL", "KFFO", "KARA", "KARG", "CWXZ", "KFFA", "KFFC", "KJDN", "KBVY", "KBVX", "KDVL", "KDVK", "KBVS", "KBVU", "KBVI", "KBVO", "KBVN", "KDVT", "KBVE", "KDVP", "CWBJ", "PAWD", "CMSI", "KGRD", "KGRF", "KGRB", "KGRI", "KGRK", "KGRR", "CWQM" ;

       Temp_instant = 273.0, 273.1, 273.2, 273.3, 273.4, 273.5,  274.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                      275.0, 273.1, 273.2, 273.3, 273.4, 273.5,  276.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                      277.0, 273.1, 273.2, 273.3, 273.4, 273.5,  278.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                      279.0, 273.1, 273.2, 273.3, 273.4, 273.5,  280.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                      281.0, 273.1, 273.2, 273.3, 273.4, 273.5,  282.0, 273.1, 273.2, 273.3, 273.4, 273.5 ;

       DewPt_instant = 273.0, 273.1, 273.2, 273.3, 273.4, 273.5,  274.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                       275.0, 273.1, 273.2, 273.3, 273.4, 273.5,  276.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                       277.0, 273.1, 273.2, 273.3, 273.4, 273.5,  278.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                       279.0, 273.1, 273.2, 273.3, 273.4, 273.5,  280.0, 273.1, 273.2, 273.3, 273.4, 273.5,
                       281.0, 273.1, 273.2, 273.3, 273.4, 273.5,  282.0, 273.1, 273.2, 273.3, 273.4, 273.5 ;

       RelHum_instant = 73.0, 73.1, 73.2, 73.3, 73.4, 73.5,  74.0, 73.1, 73.2, 73.3, 73.4, 73.5,
                        75.0, 73.1, 73.2, 73.3, 73.4, 73.5,  76.0, 73.1, 73.2, 73.3, 73.4, 73.5,
                        77.0, 73.1, 73.2, 73.3, 73.4, 73.5,  78.0, 73.1, 73.2, 73.3, 73.4, 73.5,
                        79.0, 73.1, 73.2, 73.3, 73.4, 73.5,  80.0, 73.1, 73.2, 73.3, 73.4, 73.5,
                        81.0, 73.1, 73.2, 73.3, 73.4, 73.5,  82.0, 73.1, 73.2, 73.3, 73.4, 73.5 ;
}