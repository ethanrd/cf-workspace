netcdf CF-DSG-H.4.2.1_SingleTrajectory {
dimensions:
	time = 42 ;
	name_strlen = 3 ;
variables:
	char trajectory(name_strlen) ;
		trajectory:cf_role = "trajectory_id" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1970-01-01 00:00:00" ;
	float lon(time) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(time) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	float z(time) ;
		z:standard_name = "altitude" ;
		z:long_name = "height above mean sea level" ;
		z:units = "km" ;
		z:positive = "up" ;
		z:axis = "Z" ;
	float O3(time) ;
		O3:standard_name = "mass_fraction_of_ozone_in_air" ;
		O3:long_name = "ozone concentration" ;
		O3:units = "1e-9" ;
		O3:coordinates = "time lon lat z" ;
	float NO3(time) ;
		NO3:standard_name = "mass_fraction_of_nitrate_radical_in_air" ;
		NO3:long_name = "NO3 concentration" ;
		NO3:units = "1e-9" ;
		NO3:coordinates = "time lon lat z" ;

// global attributes:
		:featureType = "trajectory" ;
		:Conventions = "CF-1.6" ;
data:

 trajectory = "AAA" ;

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42 ;

 lon = 2, 4, 6, 8, 10, 12, 14, 16, 18, 20, 22, 24, 26, 28, 30, 32, 34, 36, 
    38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 
    74, 76, 78, 80, 82, 84 ;

 lat = 3, 6, 9, 12, 15, 18, 21, 24, 27, 30, 33, 36, 39, 42, 45, 48, 51, 54, 
    57, 60, 63, 66, 69, 72, 75, 78, 81, 84, 87, 90, 93, 96, 99, 102, 105, 
    108, 111, 114, 117, 120, 123, 126 ;

 z = 4, 8, 12, 16, 20, 24, 28, 32, 36, 40, 44, 48, 52, 56, 60, 64, 68, 72, 
    76, 80, 84, 88, 92, 96, 100, 104, 108, 112, 116, 120, 124, 128, 132, 136, 
    140, 144, 148, 152, 156, 160, 164, 168 ;

 O3 = 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 65, 70, 75, 80, 85, 90, 
    95, 100, 105, 110, 115, 120, 125, 130, 135, 140, 145, 150, 155, 160, 165, 
    170, 175, 180, 185, 190, 195, 200, 205, 210 ;

 NO3 = 6, 12, 18, 24, 30, 36, 42, 48, 54, 60, 66, 72, 78, 84, 90, 96, 102, 
    108, 114, 120, 126, 132, 138, 144, 150, 156, 162, 168, 174, 180, 186, 
    192, 198, 204, 210, 216, 222, 228, 234, 240, 246, 252 ;
}
