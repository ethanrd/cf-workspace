netcdf pred_201607_test {
dimensions:
	latitude = 2584 ;
	number_of_stations = 2584 ;
	default_time_coordinate_size = 2 ;
	num_characters = 4 ;
	longitude = 2584 ;
	elev = 1 ;
	lead_times = 1 ;
	begin_end_size = 2 ;
	level = 1 ;
	plev = 1 ;
	nv = 2 ;
variables:
	int64 elev0(elev) ;
		elev0:long_name = "height above surface" ;
		elev0:units = "m" ;
		elev0:standard_name = "height" ;
		elev0:positive = "up" ;
		elev0:axis = "Z" ;
	int64 OM__phenomenonTimeInstant(lead_times, default_time_coordinate_size) ;
		OM__phenomenonTimeInstant:_FillValue = 9999LL ;
		OM__phenomenonTimeInstant:calendar = "gregorian" ;
		OM__phenomenonTimeInstant:units = "seconds since 1970-01-01 00:00:00.0" ;
		OM__phenomenonTimeInstant:standard_name = "time" ;
		OM__phenomenonTimeInstant:PROV__specializationOf = "( OM__phenomenonTime )" ;
	int64 OM__resultTime(default_time_coordinate_size) ;
		OM__resultTime:_FillValue = 9999LL ;
		OM__resultTime:calendar = "gregorian" ;
		OM__resultTime:units = "seconds since 1970-01-01 00:00:00.0" ;
		OM__resultTime:standard_name = "time" ;
		OM__resultTime:PROV__specializationOf = "( OM__resultTime )" ;
	int64 FcstRefTime(default_time_coordinate_size) ;
		FcstRefTime:_FillValue = 9999LL ;
		FcstRefTime:calendar = "gregorian" ;
		FcstRefTime:units = "seconds since 1970-01-01 00:00:00.0" ;
		FcstRefTime:standard_name = "FcstRefTime" ;
		FcstRefTime:PROV__specializationOf = "( StatPP__Data/Time/FcstRefTime )" ;
	int64 ValidTime(lead_times, default_time_coordinate_size, begin_end_size) ;
		ValidTime:_FillValue = 9999LL ;
		ValidTime:calendar = "gregorian" ;
		ValidTime:units = "seconds since 1970-01-01 00:00:00.0" ;
		ValidTime:standard_name = "time" ;
		ValidTime:PROV__specializationOf = "( StatPP__concepts/TimeBoundsSyntax/BeginEnd OM2__Data/Time/ValidTime )" ;
	int64 LeadTime(lead_times) ;
		LeadTime:_FillValue = 9999LL ;
		LeadTime:units = "seconds" ;
		LeadTime:standard_name = "forecast_period" ;
		LeadTime:PROV__specializationOf = "( StatPP__Data/Time/LeadTime )" ;
	int64 GFSModProcStep1 ;
		GFSModProcStep1:PROV__Activity = "StatPP__Methods/Ingest/DecodeGRIB2" ;
		GFSModProcStep1:long_name = "Ingest GRIB2-encoded GFS13 forecasts from NCEP repository" ;
		GFSModProcStep1:PROV__Used = "StatPP__Data/GFS13" ;
		GFSModProcStep1:units = 1LL ;
		GFSModProcStep1:standard_name = "source" ;
	int64 GFSModProcStep2 ;
		GFSModProcStep2:PROV__Activity = "StatPP__Methods/Geosp/LinInterp" ;
		GFSModProcStep2:long_name = "Apply MDL bilinear interpolation technique" ;
		GFSModProcStep2:standard_name = "source" ;
		GFSModProcStep2:units = 1LL ;
	int64 LinSmooth ;
		LinSmooth:PROV__Activity = "StatPP__Methods/LinSmooth" ;
		LinSmooth:long_name = "Linear Smoothing" ;
	int64 BiLinInterp ;
		BiLinInterp:PROV__Activity = "StatPP__Methods/InterpBiLinear" ;
		BiLinInterp:long_name = "Linear Interpolation" ;
	double Temp_instant_2_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_2_21600_3hr:_FillValue = 9999. ;
		Temp_instant_2_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_2_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_2_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_2_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_2_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_2_21600_3hr:coordinates = "elev0 station" ;
		Temp_instant_2_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_2_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_2_21600_3hr:units = "K" ;
		Temp_instant_2_21600_3hr:leadtime = 10800LL ;
	int64 plev0(plev) ;
		plev0:long_name = "pressure" ;
		plev0:units = "hPa" ;
		plev0:standard_name = "air_pressure" ;
		plev0:positive = "down" ;
		plev0:axis = "Z" ;
	double Temp_instant_1000_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_1000_21600_3hr:_FillValue = 9999. ;
		Temp_instant_1000_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_1000_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_1000_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_1000_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_1000_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_1000_21600_3hr:coordinates = "plev0 station" ;
		Temp_instant_1000_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_1000_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_1000_21600_3hr:units = "K" ;
		Temp_instant_1000_21600_3hr:leadtime = 10800LL ;
	int64 plev1(plev) ;
		plev1:long_name = "pressure" ;
		plev1:units = "hPa" ;
		plev1:standard_name = "air_pressure" ;
		plev1:positive = "down" ;
		plev1:axis = "Z" ;
	double Temp_instant_975_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_975_21600_3hr:_FillValue = 9999. ;
		Temp_instant_975_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_975_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_975_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_975_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_975_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_975_21600_3hr:coordinates = "plev1 station" ;
		Temp_instant_975_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_975_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_975_21600_3hr:units = "K" ;
		Temp_instant_975_21600_3hr:leadtime = 10800LL ;
	int64 plev2(plev) ;
		plev2:long_name = "pressure" ;
		plev2:units = "hPa" ;
		plev2:standard_name = "air_pressure" ;
		plev2:positive = "down" ;
		plev2:axis = "Z" ;
	double Temp_instant_950_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_950_21600_3hr:_FillValue = 9999. ;
		Temp_instant_950_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_950_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_950_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_950_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_950_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_950_21600_3hr:coordinates = "plev2 station" ;
		Temp_instant_950_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_950_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_950_21600_3hr:units = "K" ;
		Temp_instant_950_21600_3hr:leadtime = 10800LL ;
	int64 plev3(plev) ;
		plev3:long_name = "pressure" ;
		plev3:units = "hPa" ;
		plev3:standard_name = "air_pressure" ;
		plev3:positive = "down" ;
		plev3:axis = "Z" ;
	double Temp_instant_925_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_925_21600_3hr:_FillValue = 9999. ;
		Temp_instant_925_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_925_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_925_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_925_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_925_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_925_21600_3hr:coordinates = "plev3 station" ;
		Temp_instant_925_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_925_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_925_21600_3hr:units = "K" ;
		Temp_instant_925_21600_3hr:leadtime = 10800LL ;
	int64 plev4(plev) ;
		plev4:long_name = "pressure" ;
		plev4:units = "hPa" ;
		plev4:standard_name = "air_pressure" ;
		plev4:positive = "down" ;
		plev4:axis = "Z" ;
	double Temp_instant_850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_850_21600_3hr:_FillValue = 9999. ;
		Temp_instant_850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_850_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_850_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_850_21600_3hr:coordinates = "plev4 station" ;
		Temp_instant_850_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_850_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_850_21600_3hr:units = "K" ;
		Temp_instant_850_21600_3hr:leadtime = 10800LL ;
	int64 plev5(plev) ;
		plev5:long_name = "pressure" ;
		plev5:units = "hPa" ;
		plev5:standard_name = "air_pressure" ;
		plev5:positive = "down" ;
		plev5:axis = "Z" ;
	double Temp_instant_700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_700_21600_3hr:_FillValue = 9999. ;
		Temp_instant_700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Temp_instant_700_21600_3hr:long_name = "temperature instant" ;
		Temp_instant_700_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Temp_instant_700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Temp_instant_700_21600_3hr:coordinates = "plev5 station" ;
		Temp_instant_700_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_700_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_700_21600_3hr:units = "K" ;
		Temp_instant_700_21600_3hr:leadtime = 10800LL ;
	double DewPt_instant_2_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_2_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_2_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_2_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_2_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_2_21600_3hr:units = "K" ;
		DewPt_instant_2_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_2_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_2_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_2_21600_3hr:coordinates = "elev0 station" ;
		DewPt_instant_2_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double DewPt_instant_1000_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_1000_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_1000_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_1000_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_1000_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_1000_21600_3hr:units = "K" ;
		DewPt_instant_1000_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_1000_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_1000_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_1000_21600_3hr:coordinates = "plev0 station" ;
		DewPt_instant_1000_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double DewPt_instant_975_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_975_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_975_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_975_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_975_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_975_21600_3hr:units = "K" ;
		DewPt_instant_975_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_975_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_975_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_975_21600_3hr:coordinates = "plev1 station" ;
		DewPt_instant_975_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double DewPt_instant_950_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_950_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_950_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_950_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_950_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_950_21600_3hr:units = "K" ;
		DewPt_instant_950_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_950_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_950_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_950_21600_3hr:coordinates = "plev2 station" ;
		DewPt_instant_950_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double DewPt_instant_925_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_925_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_925_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_925_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_925_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_925_21600_3hr:units = "K" ;
		DewPt_instant_925_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_925_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_925_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_925_21600_3hr:coordinates = "plev3 station" ;
		DewPt_instant_925_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double DewPt_instant_850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_850_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_850_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_850_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_850_21600_3hr:units = "K" ;
		DewPt_instant_850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_850_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_850_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_850_21600_3hr:coordinates = "plev4 station" ;
		DewPt_instant_850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double DewPt_instant_700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		DewPt_instant_700_21600_3hr:_FillValue = 9999. ;
		DewPt_instant_700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/DewPt" ;
		DewPt_instant_700_21600_3hr:standard_name = "dew_point_temperature" ;
		DewPt_instant_700_21600_3hr:long_name = "dew point temperature" ;
		DewPt_instant_700_21600_3hr:units = "K" ;
		DewPt_instant_700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		DewPt_instant_700_21600_3hr:FcstTime_hour = 21600LL ;
		DewPt_instant_700_21600_3hr:leadtime = 10800LL ;
		DewPt_instant_700_21600_3hr:coordinates = "plev5 station" ;
		DewPt_instant_700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double RelHum_instant_2_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_2_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_2_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_2_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_2_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_2_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_2_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_2_21600_3hr:coordinates = "elev0 station" ;
		RelHum_instant_2_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_2_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_2_21600_3hr:units = "%" ;
		RelHum_instant_2_21600_3hr:leadtime = 10800LL ;
	double RelHum_instant_1000_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_1000_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_1000_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_1000_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_1000_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_1000_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_1000_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_1000_21600_3hr:coordinates = "plev0 station" ;
		RelHum_instant_1000_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_1000_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_1000_21600_3hr:units = "%" ;
		RelHum_instant_1000_21600_3hr:leadtime = 10800LL ;
	double RelHum_instant_975_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_975_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_975_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_975_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_975_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_975_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_975_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_975_21600_3hr:coordinates = "plev1 station" ;
		RelHum_instant_975_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_975_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_975_21600_3hr:units = "%" ;
		RelHum_instant_975_21600_3hr:leadtime = 10800LL ;
	double RelHum_instant_950_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_950_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_950_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_950_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_950_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_950_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_950_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_950_21600_3hr:coordinates = "plev2 station" ;
		RelHum_instant_950_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_950_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_950_21600_3hr:units = "%" ;
		RelHum_instant_950_21600_3hr:leadtime = 10800LL ;
	double RelHum_instant_925_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_925_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_925_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_925_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_925_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_925_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_925_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_925_21600_3hr:coordinates = "plev3 station" ;
		RelHum_instant_925_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_925_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_925_21600_3hr:units = "%" ;
		RelHum_instant_925_21600_3hr:leadtime = 10800LL ;
	double RelHum_instant_850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_850_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_850_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_850_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_850_21600_3hr:coordinates = "plev4 station" ;
		RelHum_instant_850_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_850_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_850_21600_3hr:units = "%" ;
		RelHum_instant_850_21600_3hr:leadtime = 10800LL ;
	double RelHum_instant_700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		RelHum_instant_700_21600_3hr:_FillValue = 9999. ;
		RelHum_instant_700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/RelHum" ;
		RelHum_instant_700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		RelHum_instant_700_21600_3hr:long_name = "relative humidity instant" ;
		RelHum_instant_700_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		RelHum_instant_700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		RelHum_instant_700_21600_3hr:coordinates = "plev5 station" ;
		RelHum_instant_700_21600_3hr:FcstTime_hour = 21600LL ;
		RelHum_instant_700_21600_3hr:standard_name = "relative_humidity" ;
		RelHum_instant_700_21600_3hr:units = "%" ;
		RelHum_instant_700_21600_3hr:leadtime = 10800LL ;
	int64 plev_bounds0(plev, nv) ;
		plev_bounds0:long_name = "pressure layer bounds" ;
		plev_bounds0:units = "hPa" ;
		plev_bounds0:standard_name = "air_pressure_layer_bounds" ;
		plev_bounds0:positive = "down" ;
		plev_bounds0:axis = "Z" ;
	int64 PressThickness ;
		PressThickness:PROV__Activity = "StatPP__Methods/Thermo/_Thick" ;
		PressThickness:long_name = "Difference of geopotential height between two isobaric levels" ;
		PressThickness:standard_name = "source" ;
		PressThickness:prototype_standard_name = "pressure_layer_thickness" ;
		PressThickness:units = "unit of observed property" ;
	double GeoHght_instant_500-700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		GeoHght_instant_500-700_21600_3hr:_FillValue = 9999. ;
		GeoHght_instant_500-700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Mass/GeoHght" ;
		GeoHght_instant_500-700_21600_3hr:FcstTime_hour = 21600LL ;
		GeoHght_instant_500-700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 PressThickness LinSmooth BiLinInterp " ;
		GeoHght_instant_500-700_21600_3hr:standard_name = "geopotential_height" ;
		GeoHght_instant_500-700_21600_3hr:coordinates = "plev_bounds0 station" ;
		GeoHght_instant_500-700_21600_3hr:long_name = "Difference of geopotential height between two isobaric levels" ;
		GeoHght_instant_500-700_21600_3hr:valid_min = 0. ;
		GeoHght_instant_500-700_21600_3hr:cell_methods = "pressure_level : PressThickness" ;
		GeoHght_instant_500-700_21600_3hr:units = "gpm" ;
		GeoHght_instant_500-700_21600_3hr:valid_max = 100000. ;
		GeoHght_instant_500-700_21600_3hr:leadtime = 10800LL ;
		GeoHght_instant_500-700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 PressThickness LinSmooth BiLinInterp )" ;
	int64 plev_bounds1(plev, nv) ;
		plev_bounds1:long_name = "pressure layer bounds" ;
		plev_bounds1:units = "hPa" ;
		plev_bounds1:standard_name = "air_pressure_layer_bounds" ;
		plev_bounds1:positive = "down" ;
		plev_bounds1:axis = "Z" ;
	double GeoHght_instant_700-850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		GeoHght_instant_700-850_21600_3hr:_FillValue = 9999. ;
		GeoHght_instant_700-850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Mass/GeoHght" ;
		GeoHght_instant_700-850_21600_3hr:FcstTime_hour = 21600LL ;
		GeoHght_instant_700-850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 PressThickness LinSmooth BiLinInterp " ;
		GeoHght_instant_700-850_21600_3hr:standard_name = "geopotential_height" ;
		GeoHght_instant_700-850_21600_3hr:coordinates = "plev_bounds1 station" ;
		GeoHght_instant_700-850_21600_3hr:long_name = "Difference of geopotential height between two isobaric levels" ;
		GeoHght_instant_700-850_21600_3hr:valid_min = 0. ;
		GeoHght_instant_700-850_21600_3hr:cell_methods = "pressure_level : PressThickness" ;
		GeoHght_instant_700-850_21600_3hr:units = "gpm" ;
		GeoHght_instant_700-850_21600_3hr:valid_max = 100000. ;
		GeoHght_instant_700-850_21600_3hr:leadtime = 10800LL ;
		GeoHght_instant_700-850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 PressThickness LinSmooth BiLinInterp )" ;
	int64 plev_bounds2(plev, nv) ;
		plev_bounds2:long_name = "pressure layer bounds" ;
		plev_bounds2:units = "hPa" ;
		plev_bounds2:standard_name = "air_pressure_layer_bounds" ;
		plev_bounds2:positive = "down" ;
		plev_bounds2:axis = "Z" ;
	double GeoHght_instant_850-1000_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		GeoHght_instant_850-1000_21600_3hr:_FillValue = 9999. ;
		GeoHght_instant_850-1000_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Mass/GeoHght" ;
		GeoHght_instant_850-1000_21600_3hr:FcstTime_hour = 21600LL ;
		GeoHght_instant_850-1000_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 PressThickness LinSmooth BiLinInterp " ;
		GeoHght_instant_850-1000_21600_3hr:standard_name = "geopotential_height" ;
		GeoHght_instant_850-1000_21600_3hr:coordinates = "plev_bounds2 station" ;
		GeoHght_instant_850-1000_21600_3hr:long_name = "Difference of geopotential height between two isobaric levels" ;
		GeoHght_instant_850-1000_21600_3hr:valid_min = 0. ;
		GeoHght_instant_850-1000_21600_3hr:cell_methods = "pressure_level : PressThickness" ;
		GeoHght_instant_850-1000_21600_3hr:units = "gpm" ;
		GeoHght_instant_850-1000_21600_3hr:valid_max = 100000. ;
		GeoHght_instant_850-1000_21600_3hr:leadtime = 10800LL ;
		GeoHght_instant_850-1000_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 PressThickness LinSmooth BiLinInterp )" ;
	int64 elev1(elev) ;
		elev1:long_name = "height above surface" ;
		elev1:units = "m" ;
		elev1:standard_name = "height" ;
		elev1:positive = "up" ;
		elev1:axis = "Z" ;
	double Uwind_instant_10_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Uwind_instant_10_21600_3hr:_FillValue = 9999. ;
		Uwind_instant_10_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/Uwind" ;
		Uwind_instant_10_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Uwind_instant_10_21600_3hr:long_name = "U wind speed instant" ;
		Uwind_instant_10_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Uwind_instant_10_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Uwind_instant_10_21600_3hr:coordinates = "elev1 station" ;
		Uwind_instant_10_21600_3hr:FcstTime_hour = 21600LL ;
		Uwind_instant_10_21600_3hr:standard_name = "eastward_wind" ;
		Uwind_instant_10_21600_3hr:units = "m s**-1" ;
		Uwind_instant_10_21600_3hr:leadtime = 10800LL ;
	double Vwind_instant_10_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Vwind_instant_10_21600_3hr:_FillValue = 9999. ;
		Vwind_instant_10_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/Vwind" ;
		Vwind_instant_10_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Vwind_instant_10_21600_3hr:long_name = "V wind speed instant" ;
		Vwind_instant_10_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Vwind_instant_10_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Vwind_instant_10_21600_3hr:coordinates = "elev1 station" ;
		Vwind_instant_10_21600_3hr:FcstTime_hour = 21600LL ;
		Vwind_instant_10_21600_3hr:standard_name = "northward_wind" ;
		Vwind_instant_10_21600_3hr:units = "m s**-1" ;
		Vwind_instant_10_21600_3hr:leadtime = 10800LL ;
	double WindSpd_instant_10_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_10_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_10_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_10_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_10_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_10_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_10_21600_3hr:valid_min = 0. ;
		WindSpd_instant_10_21600_3hr:coordinates = "elev1 station" ;
		WindSpd_instant_10_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_10_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_10_21600_3hr:units = "m/s" ;
		WindSpd_instant_10_21600_3hr:valid_max = 75. ;
		WindSpd_instant_10_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_10_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double WindSpd_instant_1000_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_1000_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_1000_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_1000_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_1000_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_1000_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_1000_21600_3hr:valid_min = 0. ;
		WindSpd_instant_1000_21600_3hr:coordinates = "plev0 station" ;
		WindSpd_instant_1000_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_1000_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_1000_21600_3hr:units = "m/s" ;
		WindSpd_instant_1000_21600_3hr:valid_max = 75. ;
		WindSpd_instant_1000_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_1000_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double WindSpd_instant_975_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_975_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_975_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_975_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_975_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_975_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_975_21600_3hr:valid_min = 0. ;
		WindSpd_instant_975_21600_3hr:coordinates = "plev1 station" ;
		WindSpd_instant_975_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_975_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_975_21600_3hr:units = "m/s" ;
		WindSpd_instant_975_21600_3hr:valid_max = 75. ;
		WindSpd_instant_975_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_975_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double WindSpd_instant_950_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_950_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_950_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_950_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_950_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_950_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_950_21600_3hr:valid_min = 0. ;
		WindSpd_instant_950_21600_3hr:coordinates = "plev2 station" ;
		WindSpd_instant_950_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_950_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_950_21600_3hr:units = "m/s" ;
		WindSpd_instant_950_21600_3hr:valid_max = 75. ;
		WindSpd_instant_950_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_950_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double WindSpd_instant_925_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_925_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_925_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_925_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_925_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_925_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_925_21600_3hr:valid_min = 0. ;
		WindSpd_instant_925_21600_3hr:coordinates = "plev3 station" ;
		WindSpd_instant_925_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_925_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_925_21600_3hr:units = "m/s" ;
		WindSpd_instant_925_21600_3hr:valid_max = 75. ;
		WindSpd_instant_925_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_925_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double WindSpd_instant_850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_850_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_850_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_850_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_850_21600_3hr:valid_min = 0. ;
		WindSpd_instant_850_21600_3hr:coordinates = "plev4 station" ;
		WindSpd_instant_850_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_850_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_850_21600_3hr:units = "m/s" ;
		WindSpd_instant_850_21600_3hr:valid_max = 75. ;
		WindSpd_instant_850_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double WindSpd_instant_700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WindSpd_instant_700_21600_3hr:_FillValue = 9999. ;
		WindSpd_instant_700_21600_3hr:comment = "Wind speed is set to -9 if winds are variable." ;
		WindSpd_instant_700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WindSpd" ;
		WindSpd_instant_700_21600_3hr:FcstTime_hour = 21600LL ;
		WindSpd_instant_700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WindSpd_instant_700_21600_3hr:valid_min = 0. ;
		WindSpd_instant_700_21600_3hr:coordinates = "plev5 station" ;
		WindSpd_instant_700_21600_3hr:long_name = "horizontal wind speed" ;
		WindSpd_instant_700_21600_3hr:standard_name = "wind_speed" ;
		WindSpd_instant_700_21600_3hr:units = "m/s" ;
		WindSpd_instant_700_21600_3hr:valid_max = 75. ;
		WindSpd_instant_700_21600_3hr:leadtime = 10800LL ;
		WindSpd_instant_700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double Wwind_instant_850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Wwind_instant_850_21600_3hr:_FillValue = 9999. ;
		Wwind_instant_850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/Wwind" ;
		Wwind_instant_850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Wwind_instant_850_21600_3hr:long_name = "vertical velocity instant" ;
		Wwind_instant_850_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Wwind_instant_850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Wwind_instant_850_21600_3hr:coordinates = "plev4 station" ;
		Wwind_instant_850_21600_3hr:FcstTime_hour = 21600LL ;
		Wwind_instant_850_21600_3hr:standard_name = "upward_air_velocity" ;
		Wwind_instant_850_21600_3hr:units = "Pa s**-1" ;
		Wwind_instant_850_21600_3hr:leadtime = 10800LL ;
	double Wwind_instant_700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Wwind_instant_700_21600_3hr:_FillValue = 9999. ;
		Wwind_instant_700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/Wwind" ;
		Wwind_instant_700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
		Wwind_instant_700_21600_3hr:long_name = "vertical velocity instant" ;
		Wwind_instant_700_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		Wwind_instant_700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		Wwind_instant_700_21600_3hr:coordinates = "plev5 station" ;
		Wwind_instant_700_21600_3hr:FcstTime_hour = 21600LL ;
		Wwind_instant_700_21600_3hr:standard_name = "upward_air_velocity" ;
		Wwind_instant_700_21600_3hr:units = "Pa s**-1" ;
		Wwind_instant_700_21600_3hr:leadtime = 10800LL ;
	int64 TempLapse ;
		TempLapse:PROV__Activity = "StatPP__Methods/Thermo/LapRate" ;
		TempLapse:long_name = "Derivative of air temperature with respect to increasing height" ;
		TempLapse:standard_name = "air_temperature_lapse_rate" ;
		TempLapse:units = "unit of observed property" ;
	double Temp_instant_500-700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_500-700_21600_3hr:_FillValue = 9999. ;
		Temp_instant_500-700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_500-700_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_500-700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 TempLapse LinSmooth BiLinInterp " ;
		Temp_instant_500-700_21600_3hr:coordinates = "plev_bounds0 station" ;
		Temp_instant_500-700_21600_3hr:long_name = "Difference in air temperature between two isobaric levels" ;
		Temp_instant_500-700_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_500-700_21600_3hr:cell_methods = "pressure_level : TempLapse" ;
		Temp_instant_500-700_21600_3hr:units = "kelvin" ;
		Temp_instant_500-700_21600_3hr:leadtime = 10800LL ;
		Temp_instant_500-700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 TempLapse LinSmooth BiLinInterp )" ;
	double Temp_instant_700-850_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_700-850_21600_3hr:_FillValue = 9999. ;
		Temp_instant_700-850_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_700-850_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_700-850_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 TempLapse LinSmooth BiLinInterp " ;
		Temp_instant_700-850_21600_3hr:coordinates = "plev_bounds1 station" ;
		Temp_instant_700-850_21600_3hr:long_name = "Difference in air temperature between two isobaric levels" ;
		Temp_instant_700-850_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_700-850_21600_3hr:cell_methods = "pressure_level : TempLapse" ;
		Temp_instant_700-850_21600_3hr:units = "kelvin" ;
		Temp_instant_700-850_21600_3hr:leadtime = 10800LL ;
		Temp_instant_700-850_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 TempLapse LinSmooth BiLinInterp )" ;
	double Temp_instant_850-1000_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		Temp_instant_850-1000_21600_3hr:_FillValue = 9999. ;
		Temp_instant_850-1000_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/Temp" ;
		Temp_instant_850-1000_21600_3hr:FcstTime_hour = 21600LL ;
		Temp_instant_850-1000_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 TempLapse LinSmooth BiLinInterp " ;
		Temp_instant_850-1000_21600_3hr:coordinates = "plev_bounds2 station" ;
		Temp_instant_850-1000_21600_3hr:long_name = "Difference in air temperature between two isobaric levels" ;
		Temp_instant_850-1000_21600_3hr:standard_name = "air_temperature" ;
		Temp_instant_850-1000_21600_3hr:cell_methods = "pressure_level : TempLapse" ;
		Temp_instant_850-1000_21600_3hr:units = "kelvin" ;
		Temp_instant_850-1000_21600_3hr:leadtime = 10800LL ;
		Temp_instant_850-1000_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 TempLapse LinSmooth BiLinInterp )" ;
	int64 elev2(elev) ;
		elev2:long_name = "height above surface" ;
		elev2:units = "m" ;
		elev2:standard_name = "height" ;
		elev2:positive = "up" ;
		elev2:axis = "Z" ;
	int64 OM__phenomenonTimePeriod3hr(lead_times, default_time_coordinate_size, begin_end_size) ;
		OM__phenomenonTimePeriod3hr:_FillValue = 9999LL ;
		OM__phenomenonTimePeriod3hr:calendar = "gregorian" ;
		OM__phenomenonTimePeriod3hr:units = "seconds since 1970-01-01 00:00:00.0" ;
		OM__phenomenonTimePeriod3hr:standard_name = "time" ;
		OM__phenomenonTimePeriod3hr:PROV__specializationOf = "( StatPP__concepts/TimeBoundsSyntax/BeginEnd OM__phenomenonTimePeriod )" ;
	int64 BoundsProcSum ;
		BoundsProcSum:PROV__Activity = "StatPP__Methods/Arith/Sum" ;
		BoundsProcSum:long_name = "summation within bounds" ;
	double TotalPrecip_sum_10800_0_21600_3hr(default_time_coordinate_size, number_of_stations) ;
		TotalPrecip_sum_10800_0_21600_3hr:_FillValue = 9999. ;
		TotalPrecip_sum_10800_0_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Wx/TotalPrecip" ;
		TotalPrecip_sum_10800_0_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 BoundsProcSum LinSmooth BiLinInterp )" ;
		TotalPrecip_sum_10800_0_21600_3hr:long_name = "total precipitation 3hr accum surface" ;
		TotalPrecip_sum_10800_0_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		TotalPrecip_sum_10800_0_21600_3hr:ancillary_variables = "OM__phenomenonTimePeriod3hr OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 BoundsProcSum LinSmooth BiLinInterp " ;
		TotalPrecip_sum_10800_0_21600_3hr:valid_min = 0. ;
		TotalPrecip_sum_10800_0_21600_3hr:coordinates = "elev2 station" ;
		TotalPrecip_sum_10800_0_21600_3hr:FcstTime_hour = 21600LL ;
		TotalPrecip_sum_10800_0_21600_3hr:standard_name = "precipitation_amount" ;
		TotalPrecip_sum_10800_0_21600_3hr:cell_methods = "default_time_coordinate_size : sum" ;
		TotalPrecip_sum_10800_0_21600_3hr:units = "kg m**-2" ;
		TotalPrecip_sum_10800_0_21600_3hr:leadtime = 10800LL ;
	double WChill_instant_2_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		WChill_instant_2_21600_3hr:_FillValue = 9999. ;
		WChill_instant_2_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moment/WChill" ;
		WChill_instant_2_21600_3hr:FcstTime_hour = 21600LL ;
		WChill_instant_2_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		WChill_instant_2_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		WChill_instant_2_21600_3hr:coordinates = "elev0 station" ;
		WChill_instant_2_21600_3hr:long_name = "wind chill" ;
		WChill_instant_2_21600_3hr:standard_name = "wind_chill_instant" ;
		WChill_instant_2_21600_3hr:units = "degF" ;
		WChill_instant_2_21600_3hr:leadtime = 10800LL ;
		WChill_instant_2_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double KIndex_instant_0_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		KIndex_instant_0_21600_3hr:_FillValue = 9999. ;
		KIndex_instant_0_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Stability/KIndex" ;
		KIndex_instant_0_21600_3hr:FcstTime_hour = 21600LL ;
		KIndex_instant_0_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		KIndex_instant_0_21600_3hr:coordinates = "elev2 station" ;
		KIndex_instant_0_21600_3hr:long_name = "atmospheric stability index K" ;
		KIndex_instant_0_21600_3hr:standard_name = "K Index" ;
		KIndex_instant_0_21600_3hr:units = "degC" ;
		KIndex_instant_0_21600_3hr:leadtime = 10800LL ;
		KIndex_instant_0_21600_3hr:OM_observedProperty = "https://codes.nws.noaa.gov/StatPP/Data/Met/Stability/KIndex" ;
		KIndex_instant_0_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double MixR_instant_700_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		MixR_instant_700_21600_3hr:_FillValue = 9999. ;
		MixR_instant_700_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Moist/MixR" ;
		MixR_instant_700_21600_3hr:FcstTime_hour = 21600LL ;
		MixR_instant_700_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		MixR_instant_700_21600_3hr:standard_name = "mixing ratio" ;
		MixR_instant_700_21600_3hr:coordinates = "plev5 station" ;
		MixR_instant_700_21600_3hr:long_name = "Mixing ratio instant" ;
		MixR_instant_700_21600_3hr:valid_min = 0. ;
		MixR_instant_700_21600_3hr:units = "g/kg" ;
		MixR_instant_700_21600_3hr:valid_max = 1000. ;
		MixR_instant_700_21600_3hr:leadtime = 10800LL ;
		MixR_instant_700_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double HtIndex_instant_2_21600_3hr(default_time_coordinate_size, number_of_stations, level) ;
		HtIndex_instant_2_21600_3hr:_FillValue = 9999. ;
		HtIndex_instant_2_21600_3hr:OM__observedProperty = "StatPP__Data/Met/Temp/HtIndex" ;
		HtIndex_instant_2_21600_3hr:FcstTime_hour = 21600LL ;
		HtIndex_instant_2_21600_3hr:filepath = "/scratch3/NCEPDEV/mdl/Emily.Schlie/inputfiles/testgfs0020160700.nc" ;
		HtIndex_instant_2_21600_3hr:ancillary_variables = "OM__phenomenonTimeInstant OM__resultTime FcstRefTime ValidTime LeadTime GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp " ;
		HtIndex_instant_2_21600_3hr:coordinates = "elev0 station" ;
		HtIndex_instant_2_21600_3hr:long_name = "heat index" ;
		HtIndex_instant_2_21600_3hr:standard_name = "heat_index" ;
		HtIndex_instant_2_21600_3hr:units = "degF" ;
		HtIndex_instant_2_21600_3hr:leadtime = 10800LL ;
		HtIndex_instant_2_21600_3hr:SOSA__usedProcedure = "( GFSModProcStep1 GFSModProcStep2 LinSmooth BiLinInterp )" ;
	double latitude(latitude) ;
		latitude:_FillValue = 9999. ;
		latitude:ancillary_variables = "" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:valid_min = -90. ;
		latitude:units = "degrees_north" ;
		latitude:valid_max = 90. ;
	double longitude(longitude) ;
		longitude:_FillValue = 9999. ;
		longitude:ancillary_variables = "" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:valid_min = -180. ;
		longitude:units = "degrees_west" ;
		longitude:valid_max = 180. ;
	char station(number_of_stations, num_characters) ;
		station:_FillValue = "_" ;
		station:comment = " Only currently archives reports from stations only if the first letter of the ICAO ID is \'K\', \'P\', \'M\', \'C\', or \'T\'. " ;
		station:ancillary_variables = "" ;
		station:long_name = "ICAO METAR call letters" ;
		station:standard_name = "platform_id" ;

// global attributes:
		:primary_variables = "Temp_instant_2_21600_3hr Temp_instant_1000_21600_3hr Temp_instant_975_21600_3hr Temp_instant_950_21600_3hr Temp_instant_925_21600_3hr Temp_instant_850_21600_3hr Temp_instant_700_21600_3hr DewPt_instant_2_21600_3hr DewPt_instant_1000_21600_3hr DewPt_instant_975_21600_3hr DewPt_instant_950_21600_3hr DewPt_instant_925_21600_3hr DewPt_instant_850_21600_3hr DewPt_instant_700_21600_3hr RelHum_instant_2_21600_3hr RelHum_instant_1000_21600_3hr RelHum_instant_975_21600_3hr RelHum_instant_950_21600_3hr RelHum_instant_925_21600_3hr RelHum_instant_850_21600_3hr RelHum_instant_700_21600_3hr GeoHght_instant_500-700_21600_3hr GeoHght_instant_700-850_21600_3hr GeoHght_instant_850-1000_21600_3hr Uwind_instant_10_21600_3hr Vwind_instant_10_21600_3hr WindSpd_instant_10_21600_3hr WindSpd_instant_1000_21600_3hr WindSpd_instant_975_21600_3hr WindSpd_instant_950_21600_3hr WindSpd_instant_925_21600_3hr WindSpd_instant_850_21600_3hr WindSpd_instant_700_21600_3hr Wwind_instant_850_21600_3hr Wwind_instant_700_21600_3hr Temp_instant_500-700_21600_3hr Temp_instant_700-850_21600_3hr Temp_instant_850-1000_21600_3hr TotalPrecip_sum_10800_0_21600_3hr WChill_instant_2_21600_3hr KIndex_instant_0_21600_3hr MixR_instant_700_21600_3hr HtIndex_instant_2_21600_3hr latitude longitude station" ;
		:version = "WISPS-1.0" ;
		:references = "" ;
		:file_id = "2e8c80c8-8e31-44fe-ba24-d231e6145a23" ;
		:url = "http://www.nws.noaa.gov/mdl/, https://sats.nws.noaa.gov/~wisps/" ;
		:organization = "NOAA/MDL/SMB" ;
		:history = "Generated on NOAA\'s Weather and Climate Operational Supercomputing System" ;
		:institution = "NOAA/National Weather Service" ;
		:Conventions = "CF-1.7 WISPS-0.2" ;

group: prefix_list {

  // group attributes:
  		:StatPP__ = "http://codes.nws.noaa.gov/StatPP/" ;
  		:OM2__ = "http://codes.nws.noaa.gov/StatPP/" ;
  		:SOSA__ = "http://www.w3.org/ns/sosa/" ;
  		:OM__ = "http://www.w3.org/ns/sosa/" ;
  		:PROV__ = "http://www.w3.org/ns/prov/#" ;
  		:StatppUncertainty__ = "http://codes.nws.noaa.gov/StatPP/Uncertainty" ;
  } // group prefix_list
}
