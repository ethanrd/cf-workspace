netcdf flag_var_byte {
  dimensions:
    obs = 1000;
  variables:
    float temp( obs );
      temp:units ="Celsius";
      temp:ancillary_variables = "temp_qc" ;
      temp:_Storage = "chunked" ;
      temp:_ChunkSizes = 100 ;
      temp:_DeflateLevel = 5 ;
      temp:_Shuffle = "true" ;
      temp:_Endianness = "little" ;
    byte temp_qc(obs);
      temp_qc:flag_values = 1b, 2b, 3b, 4b, 5b, 6b;
      temp_qc:flag_meanings = "a b c d e f";
      temp_qc:_Storage = "chunked" ;
      temp_qc:_ChunkSizes = 100 ;
      temp_qc:_DeflateLevel = 5 ;
      temp_qc:_Shuffle = "true" ;
      temp_qc:_Endianness = "little" ;

    :Conventions = "CF-1.8";

  data:
     temp =
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,            
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,            
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,            
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0,
            0.0, 5.0, 14.0, 16.0, 12.0, 18.0, 17.0, 16.0, 15.0, 14.0
             ;
     temp_qc =
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            1, 2, 3, 4, 5, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6,
            6, 6, 6, 6, 6, 6, 6, 6, 6, 6
            ;
  }
